`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/20/2024 04:29:39 PM
// Design Name: 
// Module Name: data_source
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data_source(
input aclk,
input wire m_axis_src_data_tready,
output reg [31:0] m_axis_src_data_tdata,
output reg m_axis_src_data_tvalid,
output reg m_axis_src_data_tlast,
//input tx_data_ready,
//output reg tx_data_valid,
output reg [15:0] msg_count_tx_idx,
output reg [15:0] waveform_sig_rx,
output reg [15:0] waveform_sig_loopback
    );

initial begin
msg_count_tx_idx = 0;
m_axis_src_data_tvalid = 0;
m_axis_src_data_tdata = 64'd0;
m_axis_src_data_tlast = 0;
end

always @(posedge aclk)
begin
if(m_axis_src_data_tready)
begin
m_axis_src_data_tvalid=1;
if(msg_count_tx_idx == 32768)
begin
    msg_count_tx_idx = 0;
end

case(msg_count_tx_idx)

////////////////////////////////


0: waveform_sig_loopback =-2494;
1: waveform_sig_loopback =-3133;
2: waveform_sig_loopback =-2787;
3: waveform_sig_loopback =-3483;
4: waveform_sig_loopback =-1687;
5: waveform_sig_loopback =-3578;
6: waveform_sig_loopback =-3070;
7: waveform_sig_loopback =-1822;
8: waveform_sig_loopback =-2892;
9: waveform_sig_loopback =-3382;
10: waveform_sig_loopback =-1867;
11: waveform_sig_loopback =-1953;
12: waveform_sig_loopback =-4043;
13: waveform_sig_loopback =-1672;
14: waveform_sig_loopback =-1498;
15: waveform_sig_loopback =-3694;
16: waveform_sig_loopback =-2429;
17: waveform_sig_loopback =-1235;
18: waveform_sig_loopback =-2108;
19: waveform_sig_loopback =-3640;
20: waveform_sig_loopback =-1420;
21: waveform_sig_loopback =-922;
22: waveform_sig_loopback =-3618;
23: waveform_sig_loopback =176;
24: waveform_sig_loopback =-4527;
25: waveform_sig_loopback =-2716;
26: waveform_sig_loopback =1152;
27: waveform_sig_loopback =-2636;
28: waveform_sig_loopback =-2627;
29: waveform_sig_loopback =-2359;
30: waveform_sig_loopback =-915;
31: waveform_sig_loopback =-305;
32: waveform_sig_loopback =-2852;
33: waveform_sig_loopback =-1886;
34: waveform_sig_loopback =-773;
35: waveform_sig_loopback =-1772;
36: waveform_sig_loopback =-943;
37: waveform_sig_loopback =-2291;
38: waveform_sig_loopback =-543;
39: waveform_sig_loopback =-1104;
40: waveform_sig_loopback =-1899;
41: waveform_sig_loopback =-777;
42: waveform_sig_loopback =-1175;
43: waveform_sig_loopback =-1046;
44: waveform_sig_loopback =-1649;
45: waveform_sig_loopback =211;
46: waveform_sig_loopback =-1771;
47: waveform_sig_loopback =-1347;
48: waveform_sig_loopback =254;
49: waveform_sig_loopback =-1277;
50: waveform_sig_loopback =-1520;
51: waveform_sig_loopback =374;
52: waveform_sig_loopback =-671;
53: waveform_sig_loopback =-1742;
54: waveform_sig_loopback =139;
55: waveform_sig_loopback =85;
56: waveform_sig_loopback =-1367;
57: waveform_sig_loopback =-1015;
58: waveform_sig_loopback =991;
59: waveform_sig_loopback =-290;
60: waveform_sig_loopback =-2105;
61: waveform_sig_loopback =1075;
62: waveform_sig_loopback =441;
63: waveform_sig_loopback =-1532;
64: waveform_sig_loopback =2314;
65: waveform_sig_loopback =-3295;
66: waveform_sig_loopback =-204;
67: waveform_sig_loopback =2799;
68: waveform_sig_loopback =-885;
69: waveform_sig_loopback =-609;
70: waveform_sig_loopback =-677;
71: waveform_sig_loopback =1208;
72: waveform_sig_loopback =1558;
73: waveform_sig_loopback =-1219;
74: waveform_sig_loopback =84;
75: waveform_sig_loopback =1166;
76: waveform_sig_loopback =51;
77: waveform_sig_loopback =900;
78: waveform_sig_loopback =-411;
79: waveform_sig_loopback =1158;
80: waveform_sig_loopback =859;
81: waveform_sig_loopback =121;
82: waveform_sig_loopback =889;
83: waveform_sig_loopback =875;
84: waveform_sig_loopback =530;
85: waveform_sig_loopback =469;
86: waveform_sig_loopback =2391;
87: waveform_sig_loopback =-569;
88: waveform_sig_loopback =1044;
89: waveform_sig_loopback =2120;
90: waveform_sig_loopback =341;
91: waveform_sig_loopback =786;
92: waveform_sig_loopback =1738;
93: waveform_sig_loopback =1480;
94: waveform_sig_loopback =209;
95: waveform_sig_loopback =1677;
96: waveform_sig_loopback =2338;
97: waveform_sig_loopback =239;
98: waveform_sig_loopback =972;
99: waveform_sig_loopback =2989;
100: waveform_sig_loopback =1194;
101: waveform_sig_loopback =41;
102: waveform_sig_loopback =3063;
103: waveform_sig_loopback =1921;
104: waveform_sig_loopback =656;
105: waveform_sig_loopback =4071;
106: waveform_sig_loopback =-1667;
107: waveform_sig_loopback =2116;
108: waveform_sig_loopback =4487;
109: waveform_sig_loopback =945;
110: waveform_sig_loopback =1377;
111: waveform_sig_loopback =1047;
112: waveform_sig_loopback =3155;
113: waveform_sig_loopback =3556;
114: waveform_sig_loopback =296;
115: waveform_sig_loopback =2301;
116: waveform_sig_loopback =2901;
117: waveform_sig_loopback =1769;
118: waveform_sig_loopback =3087;
119: waveform_sig_loopback =1079;
120: waveform_sig_loopback =3345;
121: waveform_sig_loopback =2755;
122: waveform_sig_loopback =1522;
123: waveform_sig_loopback =3061;
124: waveform_sig_loopback =2734;
125: waveform_sig_loopback =2213;
126: waveform_sig_loopback =2537;
127: waveform_sig_loopback =3811;
128: waveform_sig_loopback =1477;
129: waveform_sig_loopback =3144;
130: waveform_sig_loopback =3403;
131: waveform_sig_loopback =2403;
132: waveform_sig_loopback =2562;
133: waveform_sig_loopback =3574;
134: waveform_sig_loopback =3337;
135: waveform_sig_loopback =1827;
136: waveform_sig_loopback =3729;
137: waveform_sig_loopback =4101;
138: waveform_sig_loopback =1777;
139: waveform_sig_loopback =2956;
140: waveform_sig_loopback =4914;
141: waveform_sig_loopback =2661;
142: waveform_sig_loopback =1992;
143: waveform_sig_loopback =4949;
144: waveform_sig_loopback =3402;
145: waveform_sig_loopback =2845;
146: waveform_sig_loopback =5469;
147: waveform_sig_loopback =54;
148: waveform_sig_loopback =4396;
149: waveform_sig_loopback =5772;
150: waveform_sig_loopback =2846;
151: waveform_sig_loopback =3062;
152: waveform_sig_loopback =2669;
153: waveform_sig_loopback =5299;
154: waveform_sig_loopback =4876;
155: waveform_sig_loopback =2010;
156: waveform_sig_loopback =4368;
157: waveform_sig_loopback =4153;
158: waveform_sig_loopback =3767;
159: waveform_sig_loopback =4699;
160: waveform_sig_loopback =2564;
161: waveform_sig_loopback =5446;
162: waveform_sig_loopback =4001;
163: waveform_sig_loopback =3302;
164: waveform_sig_loopback =4892;
165: waveform_sig_loopback =4053;
166: waveform_sig_loopback =4004;
167: waveform_sig_loopback =4199;
168: waveform_sig_loopback =5245;
169: waveform_sig_loopback =3287;
170: waveform_sig_loopback =4676;
171: waveform_sig_loopback =4927;
172: waveform_sig_loopback =4220;
173: waveform_sig_loopback =3934;
174: waveform_sig_loopback =5304;
175: waveform_sig_loopback =4933;
176: waveform_sig_loopback =3163;
177: waveform_sig_loopback =5608;
178: waveform_sig_loopback =5560;
179: waveform_sig_loopback =3151;
180: waveform_sig_loopback =4845;
181: waveform_sig_loopback =6331;
182: waveform_sig_loopback =4092;
183: waveform_sig_loopback =3782;
184: waveform_sig_loopback =6273;
185: waveform_sig_loopback =4944;
186: waveform_sig_loopback =4533;
187: waveform_sig_loopback =6599;
188: waveform_sig_loopback =1805;
189: waveform_sig_loopback =5897;
190: waveform_sig_loopback =7054;
191: waveform_sig_loopback =4589;
192: waveform_sig_loopback =4146;
193: waveform_sig_loopback =4418;
194: waveform_sig_loopback =6818;
195: waveform_sig_loopback =5968;
196: waveform_sig_loopback =3766;
197: waveform_sig_loopback =5650;
198: waveform_sig_loopback =5481;
199: waveform_sig_loopback =5441;
200: waveform_sig_loopback =5766;
201: waveform_sig_loopback =4150;
202: waveform_sig_loopback =6927;
203: waveform_sig_loopback =5098;
204: waveform_sig_loopback =4983;
205: waveform_sig_loopback =6190;
206: waveform_sig_loopback =5336;
207: waveform_sig_loopback =5510;
208: waveform_sig_loopback =5532;
209: waveform_sig_loopback =6509;
210: waveform_sig_loopback =4769;
211: waveform_sig_loopback =5854;
212: waveform_sig_loopback =6360;
213: waveform_sig_loopback =5591;
214: waveform_sig_loopback =4991;
215: waveform_sig_loopback =7035;
216: waveform_sig_loopback =5844;
217: waveform_sig_loopback =4474;
218: waveform_sig_loopback =7214;
219: waveform_sig_loopback =6328;
220: waveform_sig_loopback =4686;
221: waveform_sig_loopback =6101;
222: waveform_sig_loopback =7278;
223: waveform_sig_loopback =5523;
224: waveform_sig_loopback =4809;
225: waveform_sig_loopback =7586;
226: waveform_sig_loopback =6131;
227: waveform_sig_loopback =5658;
228: waveform_sig_loopback =7791;
229: waveform_sig_loopback =2893;
230: waveform_sig_loopback =7122;
231: waveform_sig_loopback =8249;
232: waveform_sig_loopback =5584;
233: waveform_sig_loopback =5144;
234: waveform_sig_loopback =5866;
235: waveform_sig_loopback =7708;
236: waveform_sig_loopback =6985;
237: waveform_sig_loopback =5015;
238: waveform_sig_loopback =6542;
239: waveform_sig_loopback =6760;
240: waveform_sig_loopback =6504;
241: waveform_sig_loopback =6558;
242: waveform_sig_loopback =5559;
243: waveform_sig_loopback =7765;
244: waveform_sig_loopback =6077;
245: waveform_sig_loopback =6245;
246: waveform_sig_loopback =6887;
247: waveform_sig_loopback =6563;
248: waveform_sig_loopback =6470;
249: waveform_sig_loopback =6297;
250: waveform_sig_loopback =7771;
251: waveform_sig_loopback =5472;
252: waveform_sig_loopback =6833;
253: waveform_sig_loopback =7501;
254: waveform_sig_loopback =6109;
255: waveform_sig_loopback =6184;
256: waveform_sig_loopback =7954;
257: waveform_sig_loopback =6421;
258: waveform_sig_loopback =5681;
259: waveform_sig_loopback =8003;
260: waveform_sig_loopback =7080;
261: waveform_sig_loopback =5635;
262: waveform_sig_loopback =6908;
263: waveform_sig_loopback =8139;
264: waveform_sig_loopback =6352;
265: waveform_sig_loopback =5472;
266: waveform_sig_loopback =8568;
267: waveform_sig_loopback =6812;
268: waveform_sig_loopback =6363;
269: waveform_sig_loopback =8654;
270: waveform_sig_loopback =3461;
271: waveform_sig_loopback =8053;
272: waveform_sig_loopback =9081;
273: waveform_sig_loopback =5947;
274: waveform_sig_loopback =6059;
275: waveform_sig_loopback =6658;
276: waveform_sig_loopback =8158;
277: waveform_sig_loopback =7913;
278: waveform_sig_loopback =5433;
279: waveform_sig_loopback =7284;
280: waveform_sig_loopback =7522;
281: waveform_sig_loopback =6891;
282: waveform_sig_loopback =7326;
283: waveform_sig_loopback =6181;
284: waveform_sig_loopback =8230;
285: waveform_sig_loopback =6764;
286: waveform_sig_loopback =6787;
287: waveform_sig_loopback =7336;
288: waveform_sig_loopback =7280;
289: waveform_sig_loopback =6793;
290: waveform_sig_loopback =6941;
291: waveform_sig_loopback =8357;
292: waveform_sig_loopback =5650;
293: waveform_sig_loopback =7623;
294: waveform_sig_loopback =7890;
295: waveform_sig_loopback =6381;
296: waveform_sig_loopback =6969;
297: waveform_sig_loopback =8156;
298: waveform_sig_loopback =6842;
299: waveform_sig_loopback =6293;
300: waveform_sig_loopback =8185;
301: waveform_sig_loopback =7525;
302: waveform_sig_loopback =5996;
303: waveform_sig_loopback =7242;
304: waveform_sig_loopback =8669;
305: waveform_sig_loopback =6455;
306: waveform_sig_loopback =5857;
307: waveform_sig_loopback =9166;
308: waveform_sig_loopback =6690;
309: waveform_sig_loopback =6926;
310: waveform_sig_loopback =8956;
311: waveform_sig_loopback =3377;
312: waveform_sig_loopback =8825;
313: waveform_sig_loopback =9085;
314: waveform_sig_loopback =5989;
315: waveform_sig_loopback =6590;
316: waveform_sig_loopback =6564;
317: waveform_sig_loopback =8568;
318: waveform_sig_loopback =8115;
319: waveform_sig_loopback =5247;
320: waveform_sig_loopback =7890;
321: waveform_sig_loopback =7377;
322: waveform_sig_loopback =6996;
323: waveform_sig_loopback =7631;
324: waveform_sig_loopback =6046;
325: waveform_sig_loopback =8496;
326: waveform_sig_loopback =6797;
327: waveform_sig_loopback =6791;
328: waveform_sig_loopback =7535;
329: waveform_sig_loopback =7326;
330: waveform_sig_loopback =6651;
331: waveform_sig_loopback =7237;
332: waveform_sig_loopback =8261;
333: waveform_sig_loopback =5558;
334: waveform_sig_loopback =7941;
335: waveform_sig_loopback =7591;
336: waveform_sig_loopback =6381;
337: waveform_sig_loopback =7185;
338: waveform_sig_loopback =7753;
339: waveform_sig_loopback =7020;
340: waveform_sig_loopback =6165;
341: waveform_sig_loopback =7991;
342: waveform_sig_loopback =7770;
343: waveform_sig_loopback =5470;
344: waveform_sig_loopback =7449;
345: waveform_sig_loopback =8572;
346: waveform_sig_loopback =5940;
347: waveform_sig_loopback =6150;
348: waveform_sig_loopback =8841;
349: waveform_sig_loopback =6362;
350: waveform_sig_loopback =7093;
351: waveform_sig_loopback =8345;
352: waveform_sig_loopback =3271;
353: waveform_sig_loopback =8918;
354: waveform_sig_loopback =8470;
355: waveform_sig_loopback =5935;
356: waveform_sig_loopback =6336;
357: waveform_sig_loopback =6201;
358: waveform_sig_loopback =8602;
359: waveform_sig_loopback =7573;
360: waveform_sig_loopback =4933;
361: waveform_sig_loopback =7863;
362: waveform_sig_loopback =6709;
363: waveform_sig_loopback =6931;
364: waveform_sig_loopback =7232;
365: waveform_sig_loopback =5502;
366: waveform_sig_loopback =8402;
367: waveform_sig_loopback =6242;
368: waveform_sig_loopback =6305;
369: waveform_sig_loopback =7341;
370: waveform_sig_loopback =6667;
371: waveform_sig_loopback =6262;
372: waveform_sig_loopback =7098;
373: waveform_sig_loopback =7331;
374: waveform_sig_loopback =5362;
375: waveform_sig_loopback =7437;
376: waveform_sig_loopback =6882;
377: waveform_sig_loopback =6274;
378: waveform_sig_loopback =6271;
379: waveform_sig_loopback =7454;
380: waveform_sig_loopback =6478;
381: waveform_sig_loopback =5406;
382: waveform_sig_loopback =7769;
383: waveform_sig_loopback =6933;
384: waveform_sig_loopback =4859;
385: waveform_sig_loopback =7109;
386: waveform_sig_loopback =7773;
387: waveform_sig_loopback =5304;
388: waveform_sig_loopback =5708;
389: waveform_sig_loopback =8113;
390: waveform_sig_loopback =5609;
391: waveform_sig_loopback =6749;
392: waveform_sig_loopback =7289;
393: waveform_sig_loopback =2731;
394: waveform_sig_loopback =8464;
395: waveform_sig_loopback =7421;
396: waveform_sig_loopback =5490;
397: waveform_sig_loopback =5360;
398: waveform_sig_loopback =5532;
399: waveform_sig_loopback =8181;
400: waveform_sig_loopback =6294;
401: waveform_sig_loopback =4481;
402: waveform_sig_loopback =7117;
403: waveform_sig_loopback =5613;
404: waveform_sig_loopback =6590;
405: waveform_sig_loopback =5921;
406: waveform_sig_loopback =4924;
407: waveform_sig_loopback =7766;
408: waveform_sig_loopback =4901;
409: waveform_sig_loopback =5923;
410: waveform_sig_loopback =6272;
411: waveform_sig_loopback =5693;
412: waveform_sig_loopback =5633;
413: waveform_sig_loopback =5969;
414: waveform_sig_loopback =6470;
415: waveform_sig_loopback =4573;
416: waveform_sig_loopback =6351;
417: waveform_sig_loopback =6054;
418: waveform_sig_loopback =5175;
419: waveform_sig_loopback =5314;
420: waveform_sig_loopback =6655;
421: waveform_sig_loopback =5296;
422: waveform_sig_loopback =4363;
423: waveform_sig_loopback =6965;
424: waveform_sig_loopback =5651;
425: waveform_sig_loopback =3806;
426: waveform_sig_loopback =6321;
427: waveform_sig_loopback =6353;
428: waveform_sig_loopback =4332;
429: waveform_sig_loopback =4551;
430: waveform_sig_loopback =6913;
431: waveform_sig_loopback =4758;
432: waveform_sig_loopback =5504;
433: waveform_sig_loopback =5765;
434: waveform_sig_loopback =1980;
435: waveform_sig_loopback =7260;
436: waveform_sig_loopback =6263;
437: waveform_sig_loopback =4275;
438: waveform_sig_loopback =3822;
439: waveform_sig_loopback =5045;
440: waveform_sig_loopback =6596;
441: waveform_sig_loopback =4891;
442: waveform_sig_loopback =3672;
443: waveform_sig_loopback =5511;
444: waveform_sig_loopback =4674;
445: waveform_sig_loopback =5230;
446: waveform_sig_loopback =4426;
447: waveform_sig_loopback =4172;
448: waveform_sig_loopback =6033;
449: waveform_sig_loopback =3655;
450: waveform_sig_loopback =4868;
451: waveform_sig_loopback =4716;
452: waveform_sig_loopback =4606;
453: waveform_sig_loopback =4102;
454: waveform_sig_loopback =4777;
455: waveform_sig_loopback =5142;
456: waveform_sig_loopback =3089;
457: waveform_sig_loopback =5058;
458: waveform_sig_loopback =4736;
459: waveform_sig_loopback =3796;
460: waveform_sig_loopback =3766;
461: waveform_sig_loopback =5476;
462: waveform_sig_loopback =3658;
463: waveform_sig_loopback =3060;
464: waveform_sig_loopback =5782;
465: waveform_sig_loopback =3765;
466: waveform_sig_loopback =2792;
467: waveform_sig_loopback =4859;
468: waveform_sig_loopback =4650;
469: waveform_sig_loopback =3298;
470: waveform_sig_loopback =2871;
471: waveform_sig_loopback =5591;
472: waveform_sig_loopback =3204;
473: waveform_sig_loopback =3859;
474: waveform_sig_loopback =4769;
475: waveform_sig_loopback =119;
476: waveform_sig_loopback =5846;
477: waveform_sig_loopback =5035;
478: waveform_sig_loopback =2281;
479: waveform_sig_loopback =2776;
480: waveform_sig_loopback =3358;
481: waveform_sig_loopback =4892;
482: waveform_sig_loopback =3714;
483: waveform_sig_loopback =1790;
484: waveform_sig_loopback =4145;
485: waveform_sig_loopback =3100;
486: waveform_sig_loopback =3546;
487: waveform_sig_loopback =3014;
488: waveform_sig_loopback =2547;
489: waveform_sig_loopback =4450;
490: waveform_sig_loopback =2082;
491: waveform_sig_loopback =3250;
492: waveform_sig_loopback =3089;
493: waveform_sig_loopback =3021;
494: waveform_sig_loopback =2513;
495: waveform_sig_loopback =2932;
496: waveform_sig_loopback =3750;
497: waveform_sig_loopback =1445;
498: waveform_sig_loopback =3245;
499: waveform_sig_loopback =3345;
500: waveform_sig_loopback =1714;
501: waveform_sig_loopback =2702;
502: waveform_sig_loopback =3597;
503: waveform_sig_loopback =1549;
504: waveform_sig_loopback =2110;
505: waveform_sig_loopback =3601;
506: waveform_sig_loopback =2202;
507: waveform_sig_loopback =1250;
508: waveform_sig_loopback =2828;
509: waveform_sig_loopback =3371;
510: waveform_sig_loopback =1239;
511: waveform_sig_loopback =1280;
512: waveform_sig_loopback =4202;
513: waveform_sig_loopback =965;
514: waveform_sig_loopback =2559;
515: waveform_sig_loopback =2771;
516: waveform_sig_loopback =-1736;
517: waveform_sig_loopback =4512;
518: waveform_sig_loopback =2857;
519: waveform_sig_loopback =576;
520: waveform_sig_loopback =1143;
521: waveform_sig_loopback =1467;
522: waveform_sig_loopback =3233;
523: waveform_sig_loopback =1825;
524: waveform_sig_loopback =21;
525: waveform_sig_loopback =2406;
526: waveform_sig_loopback =1406;
527: waveform_sig_loopback =1656;
528: waveform_sig_loopback =1138;
529: waveform_sig_loopback =940;
530: waveform_sig_loopback =2321;
531: waveform_sig_loopback =563;
532: waveform_sig_loopback =1305;
533: waveform_sig_loopback =1080;
534: waveform_sig_loopback =1648;
535: waveform_sig_loopback =235;
536: waveform_sig_loopback =1535;
537: waveform_sig_loopback =1775;
538: waveform_sig_loopback =-757;
539: waveform_sig_loopback =2162;
540: waveform_sig_loopback =948;
541: waveform_sig_loopback =-88;
542: waveform_sig_loopback =1185;
543: waveform_sig_loopback =1258;
544: waveform_sig_loopback =119;
545: waveform_sig_loopback =135;
546: waveform_sig_loopback =1605;
547: waveform_sig_loopback =658;
548: waveform_sig_loopback =-988;
549: waveform_sig_loopback =1244;
550: waveform_sig_loopback =1546;
551: waveform_sig_loopback =-1051;
552: waveform_sig_loopback =-183;
553: waveform_sig_loopback =2214;
554: waveform_sig_loopback =-1120;
555: waveform_sig_loopback =1092;
556: waveform_sig_loopback =465;
557: waveform_sig_loopback =-3440;
558: waveform_sig_loopback =2884;
559: waveform_sig_loopback =697;
560: waveform_sig_loopback =-1196;
561: waveform_sig_loopback =-764;
562: waveform_sig_loopback =-502;
563: waveform_sig_loopback =1494;
564: waveform_sig_loopback =-145;
565: waveform_sig_loopback =-2136;
566: waveform_sig_loopback =789;
567: waveform_sig_loopback =-722;
568: waveform_sig_loopback =-228;
569: waveform_sig_loopback =-563;
570: waveform_sig_loopback =-1343;
571: waveform_sig_loopback =719;
572: waveform_sig_loopback =-1276;
573: waveform_sig_loopback =-979;
574: waveform_sig_loopback =-348;
575: waveform_sig_loopback =-606;
576: waveform_sig_loopback =-1745;
577: waveform_sig_loopback =135;
578: waveform_sig_loopback =-871;
579: waveform_sig_loopback =-2070;
580: waveform_sig_loopback =131;
581: waveform_sig_loopback =-1327;
582: waveform_sig_loopback =-1391;
583: waveform_sig_loopback =-1209;
584: waveform_sig_loopback =-295;
585: waveform_sig_loopback =-1851;
586: waveform_sig_loopback =-1947;
587: waveform_sig_loopback =22;
588: waveform_sig_loopback =-1503;
589: waveform_sig_loopback =-2841;
590: waveform_sig_loopback =-542;
591: waveform_sig_loopback =-357;
592: waveform_sig_loopback =-3169;
593: waveform_sig_loopback =-1829;
594: waveform_sig_loopback =243;
595: waveform_sig_loopback =-3235;
596: waveform_sig_loopback =-272;
597: waveform_sig_loopback =-2088;
598: waveform_sig_loopback =-4925;
599: waveform_sig_loopback =1250;
600: waveform_sig_loopback =-1797;
601: waveform_sig_loopback =-2589;
602: waveform_sig_loopback =-2892;
603: waveform_sig_loopback =-2307;
604: waveform_sig_loopback =-2;
605: waveform_sig_loopback =-2654;
606: waveform_sig_loopback =-3581;
607: waveform_sig_loopback =-927;
608: waveform_sig_loopback =-3005;
609: waveform_sig_loopback =-1602;
610: waveform_sig_loopback =-2695;
611: waveform_sig_loopback =-3114;
612: waveform_sig_loopback =-827;
613: waveform_sig_loopback =-3641;
614: waveform_sig_loopback =-2424;
615: waveform_sig_loopback =-2165;
616: waveform_sig_loopback =-2811;
617: waveform_sig_loopback =-3117;
618: waveform_sig_loopback =-1852;
619: waveform_sig_loopback =-2897;
620: waveform_sig_loopback =-3610;
621: waveform_sig_loopback =-1963;
622: waveform_sig_loopback =-2987;
623: waveform_sig_loopback =-3222;
624: waveform_sig_loopback =-3207;
625: waveform_sig_loopback =-1893;
626: waveform_sig_loopback =-3787;
627: waveform_sig_loopback =-3798;
628: waveform_sig_loopback =-1529;
629: waveform_sig_loopback =-3567;
630: waveform_sig_loopback =-4608;
631: waveform_sig_loopback =-2031;
632: waveform_sig_loopback =-2548;
633: waveform_sig_loopback =-4808;
634: waveform_sig_loopback =-3338;
635: waveform_sig_loopback =-1923;
636: waveform_sig_loopback =-4741;
637: waveform_sig_loopback =-1959;
638: waveform_sig_loopback =-4246;
639: waveform_sig_loopback =-6197;
640: waveform_sig_loopback =-799;
641: waveform_sig_loopback =-3487;
642: waveform_sig_loopback =-4117;
643: waveform_sig_loopback =-5134;
644: waveform_sig_loopback =-3525;
645: waveform_sig_loopback =-1866;
646: waveform_sig_loopback =-4656;
647: waveform_sig_loopback =-4789;
648: waveform_sig_loopback =-3061;
649: waveform_sig_loopback =-4554;
650: waveform_sig_loopback =-3073;
651: waveform_sig_loopback =-4890;
652: waveform_sig_loopback =-4287;
653: waveform_sig_loopback =-2712;
654: waveform_sig_loopback =-5493;
655: waveform_sig_loopback =-3665;
656: waveform_sig_loopback =-4227;
657: waveform_sig_loopback =-4297;
658: waveform_sig_loopback =-4667;
659: waveform_sig_loopback =-3797;
660: waveform_sig_loopback =-4309;
661: waveform_sig_loopback =-5223;
662: waveform_sig_loopback =-3743;
663: waveform_sig_loopback =-4356;
664: waveform_sig_loopback =-5024;
665: waveform_sig_loopback =-4744;
666: waveform_sig_loopback =-3309;
667: waveform_sig_loopback =-5718;
668: waveform_sig_loopback =-5174;
669: waveform_sig_loopback =-3009;
670: waveform_sig_loopback =-5521;
671: waveform_sig_loopback =-5819;
672: waveform_sig_loopback =-3630;
673: waveform_sig_loopback =-4367;
674: waveform_sig_loopback =-6061;
675: waveform_sig_loopback =-5070;
676: waveform_sig_loopback =-3404;
677: waveform_sig_loopback =-6097;
678: waveform_sig_loopback =-3772;
679: waveform_sig_loopback =-5710;
680: waveform_sig_loopback =-7553;
681: waveform_sig_loopback =-2504;
682: waveform_sig_loopback =-4655;
683: waveform_sig_loopback =-5990;
684: waveform_sig_loopback =-6489;
685: waveform_sig_loopback =-4591;
686: waveform_sig_loopback =-3828;
687: waveform_sig_loopback =-5889;
688: waveform_sig_loopback =-6223;
689: waveform_sig_loopback =-4718;
690: waveform_sig_loopback =-5591;
691: waveform_sig_loopback =-4798;
692: waveform_sig_loopback =-6339;
693: waveform_sig_loopback =-5337;
694: waveform_sig_loopback =-4526;
695: waveform_sig_loopback =-6632;
696: waveform_sig_loopback =-4976;
697: waveform_sig_loopback =-5843;
698: waveform_sig_loopback =-5370;
699: waveform_sig_loopback =-6214;
700: waveform_sig_loopback =-5112;
701: waveform_sig_loopback =-5493;
702: waveform_sig_loopback =-6832;
703: waveform_sig_loopback =-4975;
704: waveform_sig_loopback =-5566;
705: waveform_sig_loopback =-6682;
706: waveform_sig_loopback =-5712;
707: waveform_sig_loopback =-4770;
708: waveform_sig_loopback =-7242;
709: waveform_sig_loopback =-6046;
710: waveform_sig_loopback =-4578;
711: waveform_sig_loopback =-6830;
712: waveform_sig_loopback =-6823;
713: waveform_sig_loopback =-5060;
714: waveform_sig_loopback =-5520;
715: waveform_sig_loopback =-7251;
716: waveform_sig_loopback =-6421;
717: waveform_sig_loopback =-4368;
718: waveform_sig_loopback =-7512;
719: waveform_sig_loopback =-4937;
720: waveform_sig_loopback =-6723;
721: waveform_sig_loopback =-8856;
722: waveform_sig_loopback =-3431;
723: waveform_sig_loopback =-5789;
724: waveform_sig_loopback =-7561;
725: waveform_sig_loopback =-7051;
726: waveform_sig_loopback =-5888;
727: waveform_sig_loopback =-5094;
728: waveform_sig_loopback =-6624;
729: waveform_sig_loopback =-7666;
730: waveform_sig_loopback =-5474;
731: waveform_sig_loopback =-6658;
732: waveform_sig_loopback =-6134;
733: waveform_sig_loopback =-7025;
734: waveform_sig_loopback =-6517;
735: waveform_sig_loopback =-5660;
736: waveform_sig_loopback =-7380;
737: waveform_sig_loopback =-6261;
738: waveform_sig_loopback =-6672;
739: waveform_sig_loopback =-6310;
740: waveform_sig_loopback =-7354;
741: waveform_sig_loopback =-5814;
742: waveform_sig_loopback =-6595;
743: waveform_sig_loopback =-7777;
744: waveform_sig_loopback =-5698;
745: waveform_sig_loopback =-6544;
746: waveform_sig_loopback =-7715;
747: waveform_sig_loopback =-6231;
748: waveform_sig_loopback =-5922;
749: waveform_sig_loopback =-8082;
750: waveform_sig_loopback =-6454;
751: waveform_sig_loopback =-5907;
752: waveform_sig_loopback =-7313;
753: waveform_sig_loopback =-7676;
754: waveform_sig_loopback =-6113;
755: waveform_sig_loopback =-5827;
756: waveform_sig_loopback =-8571;
757: waveform_sig_loopback =-6833;
758: waveform_sig_loopback =-5018;
759: waveform_sig_loopback =-8749;
760: waveform_sig_loopback =-5023;
761: waveform_sig_loopback =-8040;
762: waveform_sig_loopback =-9499;
763: waveform_sig_loopback =-3673;
764: waveform_sig_loopback =-7068;
765: waveform_sig_loopback =-7958;
766: waveform_sig_loopback =-7711;
767: waveform_sig_loopback =-6817;
768: waveform_sig_loopback =-5345;
769: waveform_sig_loopback =-7596;
770: waveform_sig_loopback =-8304;
771: waveform_sig_loopback =-5897;
772: waveform_sig_loopback =-7517;
773: waveform_sig_loopback =-6624;
774: waveform_sig_loopback =-7639;
775: waveform_sig_loopback =-7232;
776: waveform_sig_loopback =-6153;
777: waveform_sig_loopback =-7934;
778: waveform_sig_loopback =-6950;
779: waveform_sig_loopback =-7274;
780: waveform_sig_loopback =-6778;
781: waveform_sig_loopback =-7988;
782: waveform_sig_loopback =-6038;
783: waveform_sig_loopback =-7605;
784: waveform_sig_loopback =-8174;
785: waveform_sig_loopback =-5626;
786: waveform_sig_loopback =-7650;
787: waveform_sig_loopback =-7912;
788: waveform_sig_loopback =-6640;
789: waveform_sig_loopback =-6578;
790: waveform_sig_loopback =-8098;
791: waveform_sig_loopback =-7377;
792: waveform_sig_loopback =-6148;
793: waveform_sig_loopback =-7477;
794: waveform_sig_loopback =-8533;
795: waveform_sig_loopback =-6014;
796: waveform_sig_loopback =-6455;
797: waveform_sig_loopback =-9042;
798: waveform_sig_loopback =-6699;
799: waveform_sig_loopback =-5847;
800: waveform_sig_loopback =-8882;
801: waveform_sig_loopback =-5026;
802: waveform_sig_loopback =-8957;
803: waveform_sig_loopback =-9295;
804: waveform_sig_loopback =-3947;
805: waveform_sig_loopback =-7603;
806: waveform_sig_loopback =-7943;
807: waveform_sig_loopback =-8202;
808: waveform_sig_loopback =-6886;
809: waveform_sig_loopback =-5371;
810: waveform_sig_loopback =-8233;
811: waveform_sig_loopback =-8257;
812: waveform_sig_loopback =-6023;
813: waveform_sig_loopback =-7923;
814: waveform_sig_loopback =-6544;
815: waveform_sig_loopback =-7919;
816: waveform_sig_loopback =-7334;
817: waveform_sig_loopback =-6104;
818: waveform_sig_loopback =-8235;
819: waveform_sig_loopback =-7046;
820: waveform_sig_loopback =-6908;
821: waveform_sig_loopback =-7328;
822: waveform_sig_loopback =-7901;
823: waveform_sig_loopback =-5854;
824: waveform_sig_loopback =-7971;
825: waveform_sig_loopback =-7647;
826: waveform_sig_loopback =-6179;
827: waveform_sig_loopback =-7670;
828: waveform_sig_loopback =-7343;
829: waveform_sig_loopback =-7119;
830: waveform_sig_loopback =-6299;
831: waveform_sig_loopback =-8044;
832: waveform_sig_loopback =-7458;
833: waveform_sig_loopback =-5602;
834: waveform_sig_loopback =-7971;
835: waveform_sig_loopback =-8160;
836: waveform_sig_loopback =-5580;
837: waveform_sig_loopback =-6839;
838: waveform_sig_loopback =-8615;
839: waveform_sig_loopback =-6508;
840: waveform_sig_loopback =-5842;
841: waveform_sig_loopback =-8523;
842: waveform_sig_loopback =-4958;
843: waveform_sig_loopback =-8871;
844: waveform_sig_loopback =-8754;
845: waveform_sig_loopback =-3818;
846: waveform_sig_loopback =-7496;
847: waveform_sig_loopback =-7466;
848: waveform_sig_loopback =-8097;
849: waveform_sig_loopback =-6549;
850: waveform_sig_loopback =-4874;
851: waveform_sig_loopback =-8330;
852: waveform_sig_loopback =-7451;
853: waveform_sig_loopback =-5869;
854: waveform_sig_loopback =-7747;
855: waveform_sig_loopback =-5685;
856: waveform_sig_loopback =-8131;
857: waveform_sig_loopback =-6523;
858: waveform_sig_loopback =-5696;
859: waveform_sig_loopback =-8250;
860: waveform_sig_loopback =-6029;
861: waveform_sig_loopback =-6826;
862: waveform_sig_loopback =-6876;
863: waveform_sig_loopback =-7089;
864: waveform_sig_loopback =-5838;
865: waveform_sig_loopback =-7175;
866: waveform_sig_loopback =-7154;
867: waveform_sig_loopback =-5904;
868: waveform_sig_loopback =-6820;
869: waveform_sig_loopback =-7091;
870: waveform_sig_loopback =-6416;
871: waveform_sig_loopback =-5777;
872: waveform_sig_loopback =-7702;
873: waveform_sig_loopback =-6665;
874: waveform_sig_loopback =-4969;
875: waveform_sig_loopback =-7657;
876: waveform_sig_loopback =-7386;
877: waveform_sig_loopback =-4783;
878: waveform_sig_loopback =-6593;
879: waveform_sig_loopback =-7708;
880: waveform_sig_loopback =-5839;
881: waveform_sig_loopback =-5400;
882: waveform_sig_loopback =-7464;
883: waveform_sig_loopback =-4576;
884: waveform_sig_loopback =-8283;
885: waveform_sig_loopback =-7635;
886: waveform_sig_loopback =-3536;
887: waveform_sig_loopback =-6448;
888: waveform_sig_loopback =-6946;
889: waveform_sig_loopback =-7459;
890: waveform_sig_loopback =-5247;
891: waveform_sig_loopback =-4629;
892: waveform_sig_loopback =-7417;
893: waveform_sig_loopback =-6406;
894: waveform_sig_loopback =-5517;
895: waveform_sig_loopback =-6447;
896: waveform_sig_loopback =-5105;
897: waveform_sig_loopback =-7441;
898: waveform_sig_loopback =-5184;
899: waveform_sig_loopback =-5405;
900: waveform_sig_loopback =-7036;
901: waveform_sig_loopback =-5113;
902: waveform_sig_loopback =-6288;
903: waveform_sig_loopback =-5609;
904: waveform_sig_loopback =-6364;
905: waveform_sig_loopback =-4906;
906: waveform_sig_loopback =-6216;
907: waveform_sig_loopback =-6272;
908: waveform_sig_loopback =-4846;
909: waveform_sig_loopback =-5786;
910: waveform_sig_loopback =-6321;
911: waveform_sig_loopback =-5255;
912: waveform_sig_loopback =-4696;
913: waveform_sig_loopback =-7024;
914: waveform_sig_loopback =-5260;
915: waveform_sig_loopback =-4085;
916: waveform_sig_loopback =-6847;
917: waveform_sig_loopback =-5859;
918: waveform_sig_loopback =-4125;
919: waveform_sig_loopback =-5463;
920: waveform_sig_loopback =-6446;
921: waveform_sig_loopback =-5087;
922: waveform_sig_loopback =-3998;
923: waveform_sig_loopback =-6546;
924: waveform_sig_loopback =-3535;
925: waveform_sig_loopback =-6933;
926: waveform_sig_loopback =-6701;
927: waveform_sig_loopback =-2208;
928: waveform_sig_loopback =-5205;
929: waveform_sig_loopback =-6256;
930: waveform_sig_loopback =-5780;
931: waveform_sig_loopback =-4213;
932: waveform_sig_loopback =-3618;
933: waveform_sig_loopback =-5895;
934: waveform_sig_loopback =-5521;
935: waveform_sig_loopback =-4098;
936: waveform_sig_loopback =-5123;
937: waveform_sig_loopback =-4216;
938: waveform_sig_loopback =-5845;
939: waveform_sig_loopback =-3988;
940: waveform_sig_loopback =-4390;
941: waveform_sig_loopback =-5453;
942: waveform_sig_loopback =-3991;
943: waveform_sig_loopback =-4928;
944: waveform_sig_loopback =-4276;
945: waveform_sig_loopback =-5111;
946: waveform_sig_loopback =-3496;
947: waveform_sig_loopback =-4819;
948: waveform_sig_loopback =-5141;
949: waveform_sig_loopback =-3351;
950: waveform_sig_loopback =-4388;
951: waveform_sig_loopback =-5293;
952: waveform_sig_loopback =-3342;
953: waveform_sig_loopback =-3784;
954: waveform_sig_loopback =-5620;
955: waveform_sig_loopback =-3414;
956: waveform_sig_loopback =-3316;
957: waveform_sig_loopback =-5017;
958: waveform_sig_loopback =-4514;
959: waveform_sig_loopback =-2875;
960: waveform_sig_loopback =-3568;
961: waveform_sig_loopback =-5548;
962: waveform_sig_loopback =-3210;
963: waveform_sig_loopback =-2529;
964: waveform_sig_loopback =-5421;
965: waveform_sig_loopback =-1583;
966: waveform_sig_loopback =-5937;
967: waveform_sig_loopback =-4908;
968: waveform_sig_loopback =-530;
969: waveform_sig_loopback =-4142;
970: waveform_sig_loopback =-4538;
971: waveform_sig_loopback =-4132;
972: waveform_sig_loopback =-2781;
973: waveform_sig_loopback =-2009;
974: waveform_sig_loopback =-4459;
975: waveform_sig_loopback =-3962;
976: waveform_sig_loopback =-2430;
977: waveform_sig_loopback =-3587;
978: waveform_sig_loopback =-2772;
979: waveform_sig_loopback =-4018;
980: waveform_sig_loopback =-2513;
981: waveform_sig_loopback =-2853;
982: waveform_sig_loopback =-3626;
983: waveform_sig_loopback =-2723;
984: waveform_sig_loopback =-3035;
985: waveform_sig_loopback =-2607;
986: waveform_sig_loopback =-3844;
987: waveform_sig_loopback =-1370;
988: waveform_sig_loopback =-3648;
989: waveform_sig_loopback =-3347;
990: waveform_sig_loopback =-1352;
991: waveform_sig_loopback =-3390;
992: waveform_sig_loopback =-3044;
993: waveform_sig_loopback =-1834;
994: waveform_sig_loopback =-2380;
995: waveform_sig_loopback =-3469;
996: waveform_sig_loopback =-2117;
997: waveform_sig_loopback =-1433;
998: waveform_sig_loopback =-3324;
999: waveform_sig_loopback =-2985;
1000: waveform_sig_loopback =-878;
1001: waveform_sig_loopback =-2125;
1002: waveform_sig_loopback =-3873;
1003: waveform_sig_loopback =-1180;
1004: waveform_sig_loopback =-1017;
1005: waveform_sig_loopback =-3644;
1006: waveform_sig_loopback =342;
1007: waveform_sig_loopback =-4615;
1008: waveform_sig_loopback =-2867;
1009: waveform_sig_loopback =1317;
1010: waveform_sig_loopback =-2790;
1011: waveform_sig_loopback =-2523;
1012: waveform_sig_loopback =-2402;
1013: waveform_sig_loopback =-1148;
1014: waveform_sig_loopback =44;
1015: waveform_sig_loopback =-3043;
1016: waveform_sig_loopback =-2035;
1017: waveform_sig_loopback =-463;
1018: waveform_sig_loopback =-2157;
1019: waveform_sig_loopback =-730;
1020: waveform_sig_loopback =-2286;
1021: waveform_sig_loopback =-890;
1022: waveform_sig_loopback =-731;
1023: waveform_sig_loopback =-2026;
1024: waveform_sig_loopback =-967;
1025: waveform_sig_loopback =-882;
1026: waveform_sig_loopback =-1300;
1027: waveform_sig_loopback =-1690;
1028: waveform_sig_loopback =520;
1029: waveform_sig_loopback =-2278;
1030: waveform_sig_loopback =-927;
1031: waveform_sig_loopback =87;
1032: waveform_sig_loopback =-1529;
1033: waveform_sig_loopback =-953;
1034: waveform_sig_loopback =-333;
1035: waveform_sig_loopback =-245;
1036: waveform_sig_loopback =-1676;
1037: waveform_sig_loopback =-351;
1038: waveform_sig_loopback =622;
1039: waveform_sig_loopback =-1642;
1040: waveform_sig_loopback =-1070;
1041: waveform_sig_loopback =1143;
1042: waveform_sig_loopback =-469;
1043: waveform_sig_loopback =-1936;
1044: waveform_sig_loopback =916;
1045: waveform_sig_loopback =444;
1046: waveform_sig_loopback =-1558;
1047: waveform_sig_loopback =2316;
1048: waveform_sig_loopback =-3229;
1049: waveform_sig_loopback =-356;
1050: waveform_sig_loopback =2989;
1051: waveform_sig_loopback =-1116;
1052: waveform_sig_loopback =-274;
1053: waveform_sig_loopback =-900;
1054: waveform_sig_loopback =1018;
1055: waveform_sig_loopback =2010;
1056: waveform_sig_loopback =-1640;
1057: waveform_sig_loopback =440;
1058: waveform_sig_loopback =1090;
1059: waveform_sig_loopback =-335;
1060: waveform_sig_loopback =1505;
1061: waveform_sig_loopback =-926;
1062: waveform_sig_loopback =1399;
1063: waveform_sig_loopback =1079;
1064: waveform_sig_loopback =-423;
1065: waveform_sig_loopback =1324;
1066: waveform_sig_loopback =687;
1067: waveform_sig_loopback =505;
1068: waveform_sig_loopback =527;
1069: waveform_sig_loopback =2071;
1070: waveform_sig_loopback =-205;
1071: waveform_sig_loopback =1061;
1072: waveform_sig_loopback =1708;
1073: waveform_sig_loopback =554;
1074: waveform_sig_loopback =916;
1075: waveform_sig_loopback =1456;
1076: waveform_sig_loopback =1753;
1077: waveform_sig_loopback =27;
1078: waveform_sig_loopback =1648;
1079: waveform_sig_loopback =2615;
1080: waveform_sig_loopback =-89;
1081: waveform_sig_loopback =1035;
1082: waveform_sig_loopback =3183;
1083: waveform_sig_loopback =1028;
1084: waveform_sig_loopback =269;
1085: waveform_sig_loopback =2874;
1086: waveform_sig_loopback =1972;
1087: waveform_sig_loopback =909;
1088: waveform_sig_loopback =3793;
1089: waveform_sig_loopback =-1386;
1090: waveform_sig_loopback =2062;
1091: waveform_sig_loopback =4224;
1092: waveform_sig_loopback =1263;
1093: waveform_sig_loopback =1359;
1094: waveform_sig_loopback =828;
1095: waveform_sig_loopback =3493;
1096: waveform_sig_loopback =3282;
1097: waveform_sig_loopback =460;
1098: waveform_sig_loopback =2484;
1099: waveform_sig_loopback =2531;
1100: waveform_sig_loopback =1991;
1101: waveform_sig_loopback =3178;
1102: waveform_sig_loopback =791;
1103: waveform_sig_loopback =3704;
1104: waveform_sig_loopback =2540;
1105: waveform_sig_loopback =1572;
1106: waveform_sig_loopback =3343;
1107: waveform_sig_loopback =2317;
1108: waveform_sig_loopback =2571;
1109: waveform_sig_loopback =2450;
1110: waveform_sig_loopback =3640;
1111: waveform_sig_loopback =1842;
1112: waveform_sig_loopback =2936;
1113: waveform_sig_loopback =3316;
1114: waveform_sig_loopback =2756;
1115: waveform_sig_loopback =2335;
1116: waveform_sig_loopback =3579;
1117: waveform_sig_loopback =3608;
1118: waveform_sig_loopback =1467;
1119: waveform_sig_loopback =3976;
1120: waveform_sig_loopback =4131;
1121: waveform_sig_loopback =1598;
1122: waveform_sig_loopback =3168;
1123: waveform_sig_loopback =4709;
1124: waveform_sig_loopback =2785;
1125: waveform_sig_loopback =2184;
1126: waveform_sig_loopback =4289;
1127: waveform_sig_loopback =3856;
1128: waveform_sig_loopback =2878;
1129: waveform_sig_loopback =5143;
1130: waveform_sig_loopback =358;
1131: waveform_sig_loopback =3893;
1132: waveform_sig_loopback =5971;
1133: waveform_sig_loopback =3183;
1134: waveform_sig_loopback =2526;
1135: waveform_sig_loopback =2821;
1136: waveform_sig_loopback =5500;
1137: waveform_sig_loopback =4451;
1138: waveform_sig_loopback =2473;
1139: waveform_sig_loopback =4031;
1140: waveform_sig_loopback =4196;
1141: waveform_sig_loopback =4039;
1142: waveform_sig_loopback =4225;
1143: waveform_sig_loopback =2911;
1144: waveform_sig_loopback =5375;
1145: waveform_sig_loopback =3843;
1146: waveform_sig_loopback =3560;
1147: waveform_sig_loopback =4760;
1148: waveform_sig_loopback =4065;
1149: waveform_sig_loopback =4234;
1150: waveform_sig_loopback =3923;
1151: waveform_sig_loopback =5342;
1152: waveform_sig_loopback =3527;
1153: waveform_sig_loopback =4272;
1154: waveform_sig_loopback =5076;
1155: waveform_sig_loopback =4379;
1156: waveform_sig_loopback =3662;
1157: waveform_sig_loopback =5526;
1158: waveform_sig_loopback =4847;
1159: waveform_sig_loopback =3076;
1160: waveform_sig_loopback =5835;
1161: waveform_sig_loopback =5192;
1162: waveform_sig_loopback =3388;
1163: waveform_sig_loopback =4886;
1164: waveform_sig_loopback =5923;
1165: waveform_sig_loopback =4579;
1166: waveform_sig_loopback =3509;
1167: waveform_sig_loopback =6113;
1168: waveform_sig_loopback =5434;
1169: waveform_sig_loopback =3973;
1170: waveform_sig_loopback =6911;
1171: waveform_sig_loopback =1990;
1172: waveform_sig_loopback =5312;
1173: waveform_sig_loopback =7513;
1174: waveform_sig_loopback =4446;
1175: waveform_sig_loopback =4043;
1176: waveform_sig_loopback =4757;
1177: waveform_sig_loopback =6401;
1178: waveform_sig_loopback =6088;
1179: waveform_sig_loopback =4123;
1180: waveform_sig_loopback =5150;
1181: waveform_sig_loopback =5865;
1182: waveform_sig_loopback =5269;
1183: waveform_sig_loopback =5625;
1184: waveform_sig_loopback =4611;
1185: waveform_sig_loopback =6385;
1186: waveform_sig_loopback =5365;
1187: waveform_sig_loopback =5149;
1188: waveform_sig_loopback =5840;
1189: waveform_sig_loopback =5583;
1190: waveform_sig_loopback =5508;
1191: waveform_sig_loopback =5289;
1192: waveform_sig_loopback =6790;
1193: waveform_sig_loopback =4580;
1194: waveform_sig_loopback =5717;
1195: waveform_sig_loopback =6591;
1196: waveform_sig_loopback =5308;
1197: waveform_sig_loopback =5106;
1198: waveform_sig_loopback =7021;
1199: waveform_sig_loopback =5677;
1200: waveform_sig_loopback =4655;
1201: waveform_sig_loopback =7111;
1202: waveform_sig_loopback =6151;
1203: waveform_sig_loopback =4987;
1204: waveform_sig_loopback =5856;
1205: waveform_sig_loopback =7195;
1206: waveform_sig_loopback =5926;
1207: waveform_sig_loopback =4399;
1208: waveform_sig_loopback =7705;
1209: waveform_sig_loopback =6277;
1210: waveform_sig_loopback =5112;
1211: waveform_sig_loopback =8423;
1212: waveform_sig_loopback =2687;
1213: waveform_sig_loopback =6734;
1214: waveform_sig_loopback =8874;
1215: waveform_sig_loopback =5022;
1216: waveform_sig_loopback =5582;
1217: waveform_sig_loopback =5769;
1218: waveform_sig_loopback =7302;
1219: waveform_sig_loopback =7607;
1220: waveform_sig_loopback =4616;
1221: waveform_sig_loopback =6620;
1222: waveform_sig_loopback =6914;
1223: waveform_sig_loopback =6109;
1224: waveform_sig_loopback =6897;
1225: waveform_sig_loopback =5491;
1226: waveform_sig_loopback =7534;
1227: waveform_sig_loopback =6336;
1228: waveform_sig_loopback =6152;
1229: waveform_sig_loopback =6725;
1230: waveform_sig_loopback =6733;
1231: waveform_sig_loopback =6389;
1232: waveform_sig_loopback =6139;
1233: waveform_sig_loopback =8055;
1234: waveform_sig_loopback =5190;
1235: waveform_sig_loopback =6947;
1236: waveform_sig_loopback =7585;
1237: waveform_sig_loopback =5793;
1238: waveform_sig_loopback =6610;
1239: waveform_sig_loopback =7593;
1240: waveform_sig_loopback =6447;
1241: waveform_sig_loopback =6033;
1242: waveform_sig_loopback =7442;
1243: waveform_sig_loopback =7475;
1244: waveform_sig_loopback =5661;
1245: waveform_sig_loopback =6526;
1246: waveform_sig_loopback =8538;
1247: waveform_sig_loopback =6149;
1248: waveform_sig_loopback =5488;
1249: waveform_sig_loopback =8738;
1250: waveform_sig_loopback =6583;
1251: waveform_sig_loopback =6446;
1252: waveform_sig_loopback =8897;
1253: waveform_sig_loopback =3242;
1254: waveform_sig_loopback =8112;
1255: waveform_sig_loopback =9072;
1256: waveform_sig_loopback =5915;
1257: waveform_sig_loopback =6391;
1258: waveform_sig_loopback =6270;
1259: waveform_sig_loopback =8278;
1260: waveform_sig_loopback =8079;
1261: waveform_sig_loopback =5198;
1262: waveform_sig_loopback =7476;
1263: waveform_sig_loopback =7445;
1264: waveform_sig_loopback =6710;
1265: waveform_sig_loopback =7612;
1266: waveform_sig_loopback =5930;
1267: waveform_sig_loopback =8160;
1268: waveform_sig_loopback =7094;
1269: waveform_sig_loopback =6453;
1270: waveform_sig_loopback =7423;
1271: waveform_sig_loopback =7405;
1272: waveform_sig_loopback =6539;
1273: waveform_sig_loopback =7233;
1274: waveform_sig_loopback =8225;
1275: waveform_sig_loopback =5516;
1276: waveform_sig_loopback =7954;
1277: waveform_sig_loopback =7481;
1278: waveform_sig_loopback =6617;
1279: waveform_sig_loopback =7026;
1280: waveform_sig_loopback =7739;
1281: waveform_sig_loopback =7390;
1282: waveform_sig_loopback =5954;
1283: waveform_sig_loopback =8030;
1284: waveform_sig_loopback =8004;
1285: waveform_sig_loopback =5634;
1286: waveform_sig_loopback =7332;
1287: waveform_sig_loopback =8773;
1288: waveform_sig_loopback =6323;
1289: waveform_sig_loopback =6151;
1290: waveform_sig_loopback =8904;
1291: waveform_sig_loopback =6738;
1292: waveform_sig_loopback =7088;
1293: waveform_sig_loopback =8829;
1294: waveform_sig_loopback =3495;
1295: waveform_sig_loopback =8740;
1296: waveform_sig_loopback =8959;
1297: waveform_sig_loopback =6315;
1298: waveform_sig_loopback =6538;
1299: waveform_sig_loopback =6356;
1300: waveform_sig_loopback =8804;
1301: waveform_sig_loopback =8097;
1302: waveform_sig_loopback =5248;
1303: waveform_sig_loopback =7965;
1304: waveform_sig_loopback =7226;
1305: waveform_sig_loopback =7078;
1306: waveform_sig_loopback =7877;
1307: waveform_sig_loopback =5692;
1308: waveform_sig_loopback =8751;
1309: waveform_sig_loopback =6859;
1310: waveform_sig_loopback =6438;
1311: waveform_sig_loopback =8001;
1312: waveform_sig_loopback =6954;
1313: waveform_sig_loopback =6825;
1314: waveform_sig_loopback =7433;
1315: waveform_sig_loopback =7751;
1316: waveform_sig_loopback =6138;
1317: waveform_sig_loopback =7638;
1318: waveform_sig_loopback =7465;
1319: waveform_sig_loopback =6877;
1320: waveform_sig_loopback =6567;
1321: waveform_sig_loopback =8087;
1322: waveform_sig_loopback =7115;
1323: waveform_sig_loopback =5774;
1324: waveform_sig_loopback =8258;
1325: waveform_sig_loopback =7566;
1326: waveform_sig_loopback =5573;
1327: waveform_sig_loopback =7346;
1328: waveform_sig_loopback =8432;
1329: waveform_sig_loopback =6042;
1330: waveform_sig_loopback =6144;
1331: waveform_sig_loopback =8629;
1332: waveform_sig_loopback =6420;
1333: waveform_sig_loopback =7176;
1334: waveform_sig_loopback =8133;
1335: waveform_sig_loopback =3474;
1336: waveform_sig_loopback =8685;
1337: waveform_sig_loopback =8352;
1338: waveform_sig_loopback =6353;
1339: waveform_sig_loopback =5849;
1340: waveform_sig_loopback =6316;
1341: waveform_sig_loopback =8812;
1342: waveform_sig_loopback =7125;
1343: waveform_sig_loopback =5416;
1344: waveform_sig_loopback =7604;
1345: waveform_sig_loopback =6627;
1346: waveform_sig_loopback =7264;
1347: waveform_sig_loopback =6878;
1348: waveform_sig_loopback =5683;
1349: waveform_sig_loopback =8510;
1350: waveform_sig_loopback =5955;
1351: waveform_sig_loopback =6633;
1352: waveform_sig_loopback =7193;
1353: waveform_sig_loopback =6555;
1354: waveform_sig_loopback =6626;
1355: waveform_sig_loopback =6629;
1356: waveform_sig_loopback =7551;
1357: waveform_sig_loopback =5604;
1358: waveform_sig_loopback =7017;
1359: waveform_sig_loopback =7125;
1360: waveform_sig_loopback =6282;
1361: waveform_sig_loopback =6072;
1362: waveform_sig_loopback =7610;
1363: waveform_sig_loopback =6434;
1364: waveform_sig_loopback =5283;
1365: waveform_sig_loopback =7911;
1366: waveform_sig_loopback =6730;
1367: waveform_sig_loopback =4982;
1368: waveform_sig_loopback =7130;
1369: waveform_sig_loopback =7397;
1370: waveform_sig_loopback =5658;
1371: waveform_sig_loopback =5600;
1372: waveform_sig_loopback =7745;
1373: waveform_sig_loopback =6148;
1374: waveform_sig_loopback =6224;
1375: waveform_sig_loopback =7468;
1376: waveform_sig_loopback =2979;
1377: waveform_sig_loopback =7706;
1378: waveform_sig_loopback =8021;
1379: waveform_sig_loopback =5340;
1380: waveform_sig_loopback =5019;
1381: waveform_sig_loopback =6029;
1382: waveform_sig_loopback =7556;
1383: waveform_sig_loopback =6557;
1384: waveform_sig_loopback =4690;
1385: waveform_sig_loopback =6551;
1386: waveform_sig_loopback =6076;
1387: waveform_sig_loopback =6330;
1388: waveform_sig_loopback =5931;
1389: waveform_sig_loopback =5135;
1390: waveform_sig_loopback =7362;
1391: waveform_sig_loopback =5128;
1392: waveform_sig_loopback =5969;
1393: waveform_sig_loopback =5982;
1394: waveform_sig_loopback =5849;
1395: waveform_sig_loopback =5671;
1396: waveform_sig_loopback =5618;
1397: waveform_sig_loopback =6773;
1398: waveform_sig_loopback =4474;
1399: waveform_sig_loopback =6065;
1400: waveform_sig_loopback =6366;
1401: waveform_sig_loopback =4961;
1402: waveform_sig_loopback =5277;
1403: waveform_sig_loopback =6759;
1404: waveform_sig_loopback =5028;
1405: waveform_sig_loopback =4633;
1406: waveform_sig_loopback =6818;
1407: waveform_sig_loopback =5473;
1408: waveform_sig_loopback =4254;
1409: waveform_sig_loopback =5923;
1410: waveform_sig_loopback =6334;
1411: waveform_sig_loopback =4796;
1412: waveform_sig_loopback =4152;
1413: waveform_sig_loopback =7077;
1414: waveform_sig_loopback =4827;
1415: waveform_sig_loopback =5086;
1416: waveform_sig_loopback =6622;
1417: waveform_sig_loopback =1474;
1418: waveform_sig_loopback =6992;
1419: waveform_sig_loopback =6922;
1420: waveform_sig_loopback =3734;
1421: waveform_sig_loopback =4221;
1422: waveform_sig_loopback =4890;
1423: waveform_sig_loopback =6334;
1424: waveform_sig_loopback =5495;
1425: waveform_sig_loopback =3241;
1426: waveform_sig_loopback =5525;
1427: waveform_sig_loopback =5022;
1428: waveform_sig_loopback =4821;
1429: waveform_sig_loopback =4830;
1430: waveform_sig_loopback =4012;
1431: waveform_sig_loopback =5940;
1432: waveform_sig_loopback =4000;
1433: waveform_sig_loopback =4643;
1434: waveform_sig_loopback =4652;
1435: waveform_sig_loopback =4780;
1436: waveform_sig_loopback =4101;
1437: waveform_sig_loopback =4393;
1438: waveform_sig_loopback =5638;
1439: waveform_sig_loopback =2844;
1440: waveform_sig_loopback =5057;
1441: waveform_sig_loopback =4955;
1442: waveform_sig_loopback =3339;
1443: waveform_sig_loopback =4454;
1444: waveform_sig_loopback =4995;
1445: waveform_sig_loopback =3659;
1446: waveform_sig_loopback =3567;
1447: waveform_sig_loopback =5081;
1448: waveform_sig_loopback =4349;
1449: waveform_sig_loopback =2701;
1450: waveform_sig_loopback =4532;
1451: waveform_sig_loopback =5148;
1452: waveform_sig_loopback =2973;
1453: waveform_sig_loopback =2977;
1454: waveform_sig_loopback =5724;
1455: waveform_sig_loopback =3046;
1456: waveform_sig_loopback =3940;
1457: waveform_sig_loopback =4967;
1458: waveform_sig_loopback =-85;
1459: waveform_sig_loopback =5841;
1460: waveform_sig_loopback =5132;
1461: waveform_sig_loopback =2253;
1462: waveform_sig_loopback =2945;
1463: waveform_sig_loopback =3138;
1464: waveform_sig_loopback =4875;
1465: waveform_sig_loopback =4050;
1466: waveform_sig_loopback =1511;
1467: waveform_sig_loopback =4251;
1468: waveform_sig_loopback =3275;
1469: waveform_sig_loopback =3236;
1470: waveform_sig_loopback =3369;
1471: waveform_sig_loopback =2250;
1472: waveform_sig_loopback =4333;
1473: waveform_sig_loopback =2608;
1474: waveform_sig_loopback =2577;
1475: waveform_sig_loopback =3258;
1476: waveform_sig_loopback =3315;
1477: waveform_sig_loopback =2168;
1478: waveform_sig_loopback =3123;
1479: waveform_sig_loopback =3486;
1480: waveform_sig_loopback =1547;
1481: waveform_sig_loopback =3633;
1482: waveform_sig_loopback =2784;
1483: waveform_sig_loopback =1966;
1484: waveform_sig_loopback =2818;
1485: waveform_sig_loopback =3284;
1486: waveform_sig_loopback =1981;
1487: waveform_sig_loopback =1779;
1488: waveform_sig_loopback =3496;
1489: waveform_sig_loopback =2673;
1490: waveform_sig_loopback =805;
1491: waveform_sig_loopback =2880;
1492: waveform_sig_loopback =3593;
1493: waveform_sig_loopback =924;
1494: waveform_sig_loopback =1424;
1495: waveform_sig_loopback =4069;
1496: waveform_sig_loopback =961;
1497: waveform_sig_loopback =2712;
1498: waveform_sig_loopback =2699;
1499: waveform_sig_loopback =-1794;
1500: waveform_sig_loopback =4615;
1501: waveform_sig_loopback =2706;
1502: waveform_sig_loopback =736;
1503: waveform_sig_loopback =1149;
1504: waveform_sig_loopback =1186;
1505: waveform_sig_loopback =3533;
1506: waveform_sig_loopback =1723;
1507: waveform_sig_loopback =-183;
1508: waveform_sig_loopback =2732;
1509: waveform_sig_loopback =1005;
1510: waveform_sig_loopback =1748;
1511: waveform_sig_loopback =1464;
1512: waveform_sig_loopback =331;
1513: waveform_sig_loopback =2810;
1514: waveform_sig_loopback =456;
1515: waveform_sig_loopback =1034;
1516: waveform_sig_loopback =1599;
1517: waveform_sig_loopback =1101;
1518: waveform_sig_loopback =487;
1519: waveform_sig_loopback =1619;
1520: waveform_sig_loopback =1414;
1521: waveform_sig_loopback =-284;
1522: waveform_sig_loopback =1778;
1523: waveform_sig_loopback =916;
1524: waveform_sig_loopback =381;
1525: waveform_sig_loopback =651;
1526: waveform_sig_loopback =1468;
1527: waveform_sig_loopback =379;
1528: waveform_sig_loopback =-293;
1529: waveform_sig_loopback =1797;
1530: waveform_sig_loopback =712;
1531: waveform_sig_loopback =-1145;
1532: waveform_sig_loopback =1372;
1533: waveform_sig_loopback =1409;
1534: waveform_sig_loopback =-1039;
1535: waveform_sig_loopback =23;
1536: waveform_sig_loopback =1859;
1537: waveform_sig_loopback =-901;
1538: waveform_sig_loopback =1126;
1539: waveform_sig_loopback =316;
1540: waveform_sig_loopback =-3252;
1541: waveform_sig_loopback =2655;
1542: waveform_sig_loopback =642;
1543: waveform_sig_loopback =-769;
1544: waveform_sig_loopback =-1157;
1545: waveform_sig_loopback =-489;
1546: waveform_sig_loopback =1812;
1547: waveform_sig_loopback =-554;
1548: waveform_sig_loopback =-1697;
1549: waveform_sig_loopback =687;
1550: waveform_sig_loopback =-973;
1551: waveform_sig_loopback =263;
1552: waveform_sig_loopback =-882;
1553: waveform_sig_loopback =-1296;
1554: waveform_sig_loopback =1017;
1555: waveform_sig_loopback =-1699;
1556: waveform_sig_loopback =-550;
1557: waveform_sig_loopback =-492;
1558: waveform_sig_loopback =-811;
1559: waveform_sig_loopback =-1283;
1560: waveform_sig_loopback =-321;
1561: waveform_sig_loopback =-649;
1562: waveform_sig_loopback =-1964;
1563: waveform_sig_loopback =-213;
1564: waveform_sig_loopback =-995;
1565: waveform_sig_loopback =-1383;
1566: waveform_sig_loopback =-1498;
1567: waveform_sig_loopback =-88;
1568: waveform_sig_loopback =-1784;
1569: waveform_sig_loopback =-2259;
1570: waveform_sig_loopback =348;
1571: waveform_sig_loopback =-1711;
1572: waveform_sig_loopback =-2806;
1573: waveform_sig_loopback =-363;
1574: waveform_sig_loopback =-854;
1575: waveform_sig_loopback =-2626;
1576: waveform_sig_loopback =-2041;
1577: waveform_sig_loopback =-78;
1578: waveform_sig_loopback =-2632;
1579: waveform_sig_loopback =-873;
1580: waveform_sig_loopback =-1708;
1581: waveform_sig_loopback =-4944;
1582: waveform_sig_loopback =720;
1583: waveform_sig_loopback =-1192;
1584: waveform_sig_loopback =-2752;
1585: waveform_sig_loopback =-3163;
1586: waveform_sig_loopback =-2006;
1587: waveform_sig_loopback =-266;
1588: waveform_sig_loopback =-2525;
1589: waveform_sig_loopback =-3313;
1590: waveform_sig_loopback =-1393;
1591: waveform_sig_loopback =-2717;
1592: waveform_sig_loopback =-1517;
1593: waveform_sig_loopback =-3010;
1594: waveform_sig_loopback =-2752;
1595: waveform_sig_loopback =-1061;
1596: waveform_sig_loopback =-3658;
1597: waveform_sig_loopback =-2094;
1598: waveform_sig_loopback =-2577;
1599: waveform_sig_loopback =-2557;
1600: waveform_sig_loopback =-3016;
1601: waveform_sig_loopback =-2300;
1602: waveform_sig_loopback =-2372;
1603: waveform_sig_loopback =-3807;
1604: waveform_sig_loopback =-2138;
1605: waveform_sig_loopback =-2561;
1606: waveform_sig_loopback =-3519;
1607: waveform_sig_loopback =-3151;
1608: waveform_sig_loopback =-1722;
1609: waveform_sig_loopback =-3991;
1610: waveform_sig_loopback =-3693;
1611: waveform_sig_loopback =-1504;
1612: waveform_sig_loopback =-3727;
1613: waveform_sig_loopback =-4287;
1614: waveform_sig_loopback =-2258;
1615: waveform_sig_loopback =-2676;
1616: waveform_sig_loopback =-4301;
1617: waveform_sig_loopback =-3909;
1618: waveform_sig_loopback =-1732;
1619: waveform_sig_loopback =-4445;
1620: waveform_sig_loopback =-2688;
1621: waveform_sig_loopback =-3448;
1622: waveform_sig_loopback =-6632;
1623: waveform_sig_loopback =-1070;
1624: waveform_sig_loopback =-2827;
1625: waveform_sig_loopback =-4675;
1626: waveform_sig_loopback =-4832;
1627: waveform_sig_loopback =-3464;
1628: waveform_sig_loopback =-2331;
1629: waveform_sig_loopback =-4027;
1630: waveform_sig_loopback =-5042;
1631: waveform_sig_loopback =-3239;
1632: waveform_sig_loopback =-4045;
1633: waveform_sig_loopback =-3542;
1634: waveform_sig_loopback =-4593;
1635: waveform_sig_loopback =-4227;
1636: waveform_sig_loopback =-3106;
1637: waveform_sig_loopback =-5032;
1638: waveform_sig_loopback =-3771;
1639: waveform_sig_loopback =-4327;
1640: waveform_sig_loopback =-4041;
1641: waveform_sig_loopback =-4838;
1642: waveform_sig_loopback =-3826;
1643: waveform_sig_loopback =-3976;
1644: waveform_sig_loopback =-5550;
1645: waveform_sig_loopback =-3649;
1646: waveform_sig_loopback =-4092;
1647: waveform_sig_loopback =-5401;
1648: waveform_sig_loopback =-4462;
1649: waveform_sig_loopback =-3359;
1650: waveform_sig_loopback =-5881;
1651: waveform_sig_loopback =-4797;
1652: waveform_sig_loopback =-3400;
1653: waveform_sig_loopback =-5326;
1654: waveform_sig_loopback =-5595;
1655: waveform_sig_loopback =-4173;
1656: waveform_sig_loopback =-3881;
1657: waveform_sig_loopback =-6077;
1658: waveform_sig_loopback =-5486;
1659: waveform_sig_loopback =-2826;
1660: waveform_sig_loopback =-6444;
1661: waveform_sig_loopback =-3824;
1662: waveform_sig_loopback =-5087;
1663: waveform_sig_loopback =-8279;
1664: waveform_sig_loopback =-2123;
1665: waveform_sig_loopback =-4630;
1666: waveform_sig_loopback =-6319;
1667: waveform_sig_loopback =-5940;
1668: waveform_sig_loopback =-5112;
1669: waveform_sig_loopback =-3774;
1670: waveform_sig_loopback =-5479;
1671: waveform_sig_loopback =-6733;
1672: waveform_sig_loopback =-4405;
1673: waveform_sig_loopback =-5575;
1674: waveform_sig_loopback =-5139;
1675: waveform_sig_loopback =-5784;
1676: waveform_sig_loopback =-5691;
1677: waveform_sig_loopback =-4532;
1678: waveform_sig_loopback =-6283;
1679: waveform_sig_loopback =-5407;
1680: waveform_sig_loopback =-5616;
1681: waveform_sig_loopback =-5256;
1682: waveform_sig_loopback =-6495;
1683: waveform_sig_loopback =-4907;
1684: waveform_sig_loopback =-5440;
1685: waveform_sig_loopback =-7092;
1686: waveform_sig_loopback =-4643;
1687: waveform_sig_loopback =-5742;
1688: waveform_sig_loopback =-6735;
1689: waveform_sig_loopback =-5403;
1690: waveform_sig_loopback =-5142;
1691: waveform_sig_loopback =-6930;
1692: waveform_sig_loopback =-5965;
1693: waveform_sig_loopback =-5018;
1694: waveform_sig_loopback =-6186;
1695: waveform_sig_loopback =-7153;
1696: waveform_sig_loopback =-5276;
1697: waveform_sig_loopback =-4843;
1698: waveform_sig_loopback =-7834;
1699: waveform_sig_loopback =-6172;
1700: waveform_sig_loopback =-4213;
1701: waveform_sig_loopback =-7943;
1702: waveform_sig_loopback =-4454;
1703: waveform_sig_loopback =-6923;
1704: waveform_sig_loopback =-9085;
1705: waveform_sig_loopback =-3086;
1706: waveform_sig_loopback =-6194;
1707: waveform_sig_loopback =-7153;
1708: waveform_sig_loopback =-7186;
1709: waveform_sig_loopback =-6251;
1710: waveform_sig_loopback =-4644;
1711: waveform_sig_loopback =-6777;
1712: waveform_sig_loopback =-7787;
1713: waveform_sig_loopback =-5319;
1714: waveform_sig_loopback =-6775;
1715: waveform_sig_loopback =-6189;
1716: waveform_sig_loopback =-6812;
1717: waveform_sig_loopback =-6873;
1718: waveform_sig_loopback =-5474;
1719: waveform_sig_loopback =-7181;
1720: waveform_sig_loopback =-6715;
1721: waveform_sig_loopback =-6290;
1722: waveform_sig_loopback =-6416;
1723: waveform_sig_loopback =-7643;
1724: waveform_sig_loopback =-5328;
1725: waveform_sig_loopback =-7041;
1726: waveform_sig_loopback =-7660;
1727: waveform_sig_loopback =-5368;
1728: waveform_sig_loopback =-7205;
1729: waveform_sig_loopback =-7049;
1730: waveform_sig_loopback =-6702;
1731: waveform_sig_loopback =-5973;
1732: waveform_sig_loopback =-7493;
1733: waveform_sig_loopback =-7317;
1734: waveform_sig_loopback =-5432;
1735: waveform_sig_loopback =-7238;
1736: waveform_sig_loopback =-8175;
1737: waveform_sig_loopback =-5685;
1738: waveform_sig_loopback =-6092;
1739: waveform_sig_loopback =-8524;
1740: waveform_sig_loopback =-6769;
1741: waveform_sig_loopback =-5227;
1742: waveform_sig_loopback =-8592;
1743: waveform_sig_loopback =-5089;
1744: waveform_sig_loopback =-8020;
1745: waveform_sig_loopback =-9598;
1746: waveform_sig_loopback =-3719;
1747: waveform_sig_loopback =-7168;
1748: waveform_sig_loopback =-7687;
1749: waveform_sig_loopback =-7958;
1750: waveform_sig_loopback =-7030;
1751: waveform_sig_loopback =-4965;
1752: waveform_sig_loopback =-7874;
1753: waveform_sig_loopback =-8343;
1754: waveform_sig_loopback =-5672;
1755: waveform_sig_loopback =-7893;
1756: waveform_sig_loopback =-6266;
1757: waveform_sig_loopback =-7725;
1758: waveform_sig_loopback =-7560;
1759: waveform_sig_loopback =-5605;
1760: waveform_sig_loopback =-8407;
1761: waveform_sig_loopback =-6833;
1762: waveform_sig_loopback =-6775;
1763: waveform_sig_loopback =-7393;
1764: waveform_sig_loopback =-7591;
1765: waveform_sig_loopback =-6190;
1766: waveform_sig_loopback =-7609;
1767: waveform_sig_loopback =-7687;
1768: waveform_sig_loopback =-6375;
1769: waveform_sig_loopback =-7337;
1770: waveform_sig_loopback =-7583;
1771: waveform_sig_loopback =-7165;
1772: waveform_sig_loopback =-6152;
1773: waveform_sig_loopback =-8240;
1774: waveform_sig_loopback =-7567;
1775: waveform_sig_loopback =-5661;
1776: waveform_sig_loopback =-7859;
1777: waveform_sig_loopback =-8383;
1778: waveform_sig_loopback =-5860;
1779: waveform_sig_loopback =-6676;
1780: waveform_sig_loopback =-8795;
1781: waveform_sig_loopback =-6838;
1782: waveform_sig_loopback =-5832;
1783: waveform_sig_loopback =-8676;
1784: waveform_sig_loopback =-5272;
1785: waveform_sig_loopback =-8745;
1786: waveform_sig_loopback =-9230;
1787: waveform_sig_loopback =-4206;
1788: waveform_sig_loopback =-7531;
1789: waveform_sig_loopback =-7610;
1790: waveform_sig_loopback =-8559;
1791: waveform_sig_loopback =-6705;
1792: waveform_sig_loopback =-5268;
1793: waveform_sig_loopback =-8438;
1794: waveform_sig_loopback =-7776;
1795: waveform_sig_loopback =-6331;
1796: waveform_sig_loopback =-7906;
1797: waveform_sig_loopback =-6133;
1798: waveform_sig_loopback =-8375;
1799: waveform_sig_loopback =-6973;
1800: waveform_sig_loopback =-6027;
1801: waveform_sig_loopback =-8602;
1802: waveform_sig_loopback =-6410;
1803: waveform_sig_loopback =-7364;
1804: waveform_sig_loopback =-7183;
1805: waveform_sig_loopback =-7572;
1806: waveform_sig_loopback =-6418;
1807: waveform_sig_loopback =-7333;
1808: waveform_sig_loopback =-7891;
1809: waveform_sig_loopback =-6294;
1810: waveform_sig_loopback =-7204;
1811: waveform_sig_loopback =-7679;
1812: waveform_sig_loopback =-7003;
1813: waveform_sig_loopback =-6119;
1814: waveform_sig_loopback =-8198;
1815: waveform_sig_loopback =-7385;
1816: waveform_sig_loopback =-5461;
1817: waveform_sig_loopback =-8091;
1818: waveform_sig_loopback =-8073;
1819: waveform_sig_loopback =-5573;
1820: waveform_sig_loopback =-6971;
1821: waveform_sig_loopback =-8306;
1822: waveform_sig_loopback =-7001;
1823: waveform_sig_loopback =-5703;
1824: waveform_sig_loopback =-8091;
1825: waveform_sig_loopback =-5594;
1826: waveform_sig_loopback =-8573;
1827: waveform_sig_loopback =-8769;
1828: waveform_sig_loopback =-4189;
1829: waveform_sig_loopback =-6896;
1830: waveform_sig_loopback =-7965;
1831: waveform_sig_loopback =-8171;
1832: waveform_sig_loopback =-5930;
1833: waveform_sig_loopback =-5674;
1834: waveform_sig_loopback =-7788;
1835: waveform_sig_loopback =-7577;
1836: waveform_sig_loopback =-6202;
1837: waveform_sig_loopback =-7133;
1838: waveform_sig_loopback =-6314;
1839: waveform_sig_loopback =-7816;
1840: waveform_sig_loopback =-6372;
1841: waveform_sig_loopback =-6087;
1842: waveform_sig_loopback =-7921;
1843: waveform_sig_loopback =-6127;
1844: waveform_sig_loopback =-6914;
1845: waveform_sig_loopback =-6654;
1846: waveform_sig_loopback =-7255;
1847: waveform_sig_loopback =-5897;
1848: waveform_sig_loopback =-6862;
1849: waveform_sig_loopback =-7454;
1850: waveform_sig_loopback =-5915;
1851: waveform_sig_loopback =-6446;
1852: waveform_sig_loopback =-7481;
1853: waveform_sig_loopback =-6292;
1854: waveform_sig_loopback =-5597;
1855: waveform_sig_loopback =-8059;
1856: waveform_sig_loopback =-6281;
1857: waveform_sig_loopback =-5292;
1858: waveform_sig_loopback =-7567;
1859: waveform_sig_loopback =-7067;
1860: waveform_sig_loopback =-5404;
1861: waveform_sig_loopback =-6083;
1862: waveform_sig_loopback =-7743;
1863: waveform_sig_loopback =-6318;
1864: waveform_sig_loopback =-4807;
1865: waveform_sig_loopback =-7821;
1866: waveform_sig_loopback =-4676;
1867: waveform_sig_loopback =-7678;
1868: waveform_sig_loopback =-8283;
1869: waveform_sig_loopback =-3285;
1870: waveform_sig_loopback =-6279;
1871: waveform_sig_loopback =-7403;
1872: waveform_sig_loopback =-6919;
1873: waveform_sig_loopback =-5614;
1874: waveform_sig_loopback =-4802;
1875: waveform_sig_loopback =-6824;
1876: waveform_sig_loopback =-7033;
1877: waveform_sig_loopback =-5184;
1878: waveform_sig_loopback =-6425;
1879: waveform_sig_loopback =-5537;
1880: waveform_sig_loopback =-6827;
1881: waveform_sig_loopback =-5667;
1882: waveform_sig_loopback =-5324;
1883: waveform_sig_loopback =-6816;
1884: waveform_sig_loopback =-5426;
1885: waveform_sig_loopback =-6074;
1886: waveform_sig_loopback =-5625;
1887: waveform_sig_loopback =-6550;
1888: waveform_sig_loopback =-4828;
1889: waveform_sig_loopback =-5992;
1890: waveform_sig_loopback =-6698;
1891: waveform_sig_loopback =-4578;
1892: waveform_sig_loopback =-5796;
1893: waveform_sig_loopback =-6590;
1894: waveform_sig_loopback =-4857;
1895: waveform_sig_loopback =-5104;
1896: waveform_sig_loopback =-6759;
1897: waveform_sig_loopback =-5177;
1898: waveform_sig_loopback =-4589;
1899: waveform_sig_loopback =-6179;
1900: waveform_sig_loopback =-6283;
1901: waveform_sig_loopback =-4277;
1902: waveform_sig_loopback =-4882;
1903: waveform_sig_loopback =-6965;
1904: waveform_sig_loopback =-4890;
1905: waveform_sig_loopback =-3793;
1906: waveform_sig_loopback =-6934;
1907: waveform_sig_loopback =-3142;
1908: waveform_sig_loopback =-6987;
1909: waveform_sig_loopback =-7029;
1910: waveform_sig_loopback =-1810;
1911: waveform_sig_loopback =-5588;
1912: waveform_sig_loopback =-6032;
1913: waveform_sig_loopback =-5633;
1914: waveform_sig_loopback =-4691;
1915: waveform_sig_loopback =-3279;
1916: waveform_sig_loopback =-5886;
1917: waveform_sig_loopback =-5797;
1918: waveform_sig_loopback =-3746;
1919: waveform_sig_loopback =-5448;
1920: waveform_sig_loopback =-4169;
1921: waveform_sig_loopback =-5572;
1922: waveform_sig_loopback =-4485;
1923: waveform_sig_loopback =-3994;
1924: waveform_sig_loopback =-5525;
1925: waveform_sig_loopback =-4318;
1926: waveform_sig_loopback =-4536;
1927: waveform_sig_loopback =-4392;
1928: waveform_sig_loopback =-5410;
1929: waveform_sig_loopback =-3106;
1930: waveform_sig_loopback =-5054;
1931: waveform_sig_loopback =-5147;
1932: waveform_sig_loopback =-3060;
1933: waveform_sig_loopback =-4864;
1934: waveform_sig_loopback =-4763;
1935: waveform_sig_loopback =-3723;
1936: waveform_sig_loopback =-3884;
1937: waveform_sig_loopback =-4986;
1938: waveform_sig_loopback =-4129;
1939: waveform_sig_loopback =-2995;
1940: waveform_sig_loopback =-4800;
1941: waveform_sig_loopback =-4989;
1942: waveform_sig_loopback =-2516;
1943: waveform_sig_loopback =-3727;
1944: waveform_sig_loopback =-5583;
1945: waveform_sig_loopback =-3084;
1946: waveform_sig_loopback =-2708;
1947: waveform_sig_loopback =-5379;
1948: waveform_sig_loopback =-1456;
1949: waveform_sig_loopback =-6066;
1950: waveform_sig_loopback =-5003;
1951: waveform_sig_loopback =-323;
1952: waveform_sig_loopback =-4446;
1953: waveform_sig_loopback =-4181;
1954: waveform_sig_loopback =-4357;
1955: waveform_sig_loopback =-3069;
1956: waveform_sig_loopback =-1494;
1957: waveform_sig_loopback =-4882;
1958: waveform_sig_loopback =-3832;
1959: waveform_sig_loopback =-2271;
1960: waveform_sig_loopback =-4094;
1961: waveform_sig_loopback =-2211;
1962: waveform_sig_loopback =-4326;
1963: waveform_sig_loopback =-2718;
1964: waveform_sig_loopback =-2296;
1965: waveform_sig_loopback =-4127;
1966: waveform_sig_loopback =-2536;
1967: waveform_sig_loopback =-2888;
1968: waveform_sig_loopback =-2988;
1969: waveform_sig_loopback =-3550;
1970: waveform_sig_loopback =-1511;
1971: waveform_sig_loopback =-3684;
1972: waveform_sig_loopback =-3093;
1973: waveform_sig_loopback =-1685;
1974: waveform_sig_loopback =-3236;
1975: waveform_sig_loopback =-2815;
1976: waveform_sig_loopback =-2339;
1977: waveform_sig_loopback =-1992;
1978: waveform_sig_loopback =-3367;
1979: waveform_sig_loopback =-2611;
1980: waveform_sig_loopback =-929;
1981: waveform_sig_loopback =-3469;
1982: waveform_sig_loopback =-3173;
1983: waveform_sig_loopback =-522;
1984: waveform_sig_loopback =-2515;
1985: waveform_sig_loopback =-3523;
1986: waveform_sig_loopback =-1277;
1987: waveform_sig_loopback =-1354;
1988: waveform_sig_loopback =-3198;
1989: waveform_sig_loopback =60;
1990: waveform_sig_loopback =-4493;
1991: waveform_sig_loopback =-2797;
1992: waveform_sig_loopback =1063;
1993: waveform_sig_loopback =-2538;
1994: waveform_sig_loopback =-2418;
1995: waveform_sig_loopback =-2791;
1996: waveform_sig_loopback =-900;
1997: waveform_sig_loopback =46;
1998: waveform_sig_loopback =-3235;
1999: waveform_sig_loopback =-1671;
2000: waveform_sig_loopback =-794;
2001: waveform_sig_loopback =-2152;
2002: waveform_sig_loopback =-295;
2003: waveform_sig_loopback =-2822;
2004: waveform_sig_loopback =-645;
2005: waveform_sig_loopback =-605;
2006: waveform_sig_loopback =-2442;
2007: waveform_sig_loopback =-454;
2008: waveform_sig_loopback =-1268;
2009: waveform_sig_loopback =-1267;
2010: waveform_sig_loopback =-1374;
2011: waveform_sig_loopback =-44;
2012: waveform_sig_loopback =-1781;
2013: waveform_sig_loopback =-1062;
2014: waveform_sig_loopback =-264;
2015: waveform_sig_loopback =-976;
2016: waveform_sig_loopback =-1293;
2017: waveform_sig_loopback =-485;
2018: waveform_sig_loopback =188;
2019: waveform_sig_loopback =-2028;
2020: waveform_sig_loopback =-328;
2021: waveform_sig_loopback =800;
2022: waveform_sig_loopback =-1863;
2023: waveform_sig_loopback =-906;
2024: waveform_sig_loopback =1069;
2025: waveform_sig_loopback =-658;
2026: waveform_sig_loopback =-1546;
2027: waveform_sig_loopback =511;
2028: waveform_sig_loopback =476;
2029: waveform_sig_loopback =-1175;
2030: waveform_sig_loopback =1774;
2031: waveform_sig_loopback =-2659;
2032: waveform_sig_loopback =-673;
2033: waveform_sig_loopback =2707;
2034: waveform_sig_loopback =-477;
2035: waveform_sig_loopback =-675;
2036: waveform_sig_loopback =-942;
2037: waveform_sig_loopback =1263;
2038: waveform_sig_loopback =1588;
2039: waveform_sig_loopback =-1240;
2040: waveform_sig_loopback =351;
2041: waveform_sig_loopback =739;
2042: waveform_sig_loopback =110;
2043: waveform_sig_loopback =1400;
2044: waveform_sig_loopback =-1074;
2045: waveform_sig_loopback =1690;
2046: waveform_sig_loopback =821;
2047: waveform_sig_loopback =-295;
2048: waveform_sig_loopback =1460;
2049: waveform_sig_loopback =391;
2050: waveform_sig_loopback =954;
2051: waveform_sig_loopback =342;
2052: waveform_sig_loopback =1811;
2053: waveform_sig_loopback =349;
2054: waveform_sig_loopback =597;
2055: waveform_sig_loopback =1766;
2056: waveform_sig_loopback =976;
2057: waveform_sig_loopback =308;
2058: waveform_sig_loopback =1836;
2059: waveform_sig_loopback =1778;
2060: waveform_sig_loopback =-213;
2061: waveform_sig_loopback =1950;
2062: waveform_sig_loopback =2313;
2063: waveform_sig_loopback =130;
2064: waveform_sig_loopback =1142;
2065: waveform_sig_loopback =2763;
2066: waveform_sig_loopback =1381;
2067: waveform_sig_loopback =279;
2068: waveform_sig_loopback =2439;
2069: waveform_sig_loopback =2403;
2070: waveform_sig_loopback =618;
2071: waveform_sig_loopback =3649;
2072: waveform_sig_loopback =-846;
2073: waveform_sig_loopback =1349;
2074: waveform_sig_loopback =4452;
2075: waveform_sig_loopback =1515;
2076: waveform_sig_loopback =849;
2077: waveform_sig_loopback =1209;
2078: waveform_sig_loopback =3233;
2079: waveform_sig_loopback =3078;
2080: waveform_sig_loopback =1016;
2081: waveform_sig_loopback =1892;
2082: waveform_sig_loopback =2713;
2083: waveform_sig_loopback =2177;
2084: waveform_sig_loopback =2676;
2085: waveform_sig_loopback =1272;
2086: waveform_sig_loopback =3345;
2087: waveform_sig_loopback =2429;
2088: waveform_sig_loopback =1934;
2089: waveform_sig_loopback =2911;
2090: waveform_sig_loopback =2420;
2091: waveform_sig_loopback =2796;
2092: waveform_sig_loopback =1992;
2093: waveform_sig_loopback =3935;
2094: waveform_sig_loopback =1866;
2095: waveform_sig_loopback =2503;
2096: waveform_sig_loopback =3731;
2097: waveform_sig_loopback =2562;
2098: waveform_sig_loopback =2202;
2099: waveform_sig_loopback =3758;
2100: waveform_sig_loopback =3416;
2101: waveform_sig_loopback =1576;
2102: waveform_sig_loopback =3949;
2103: waveform_sig_loopback =3860;
2104: waveform_sig_loopback =1988;
2105: waveform_sig_loopback =3112;
2106: waveform_sig_loopback =4264;
2107: waveform_sig_loopback =3393;
2108: waveform_sig_loopback =1854;
2109: waveform_sig_loopback =4276;
2110: waveform_sig_loopback =4372;
2111: waveform_sig_loopback =2037;
2112: waveform_sig_loopback =5786;
2113: waveform_sig_loopback =613;
2114: waveform_sig_loopback =3153;
2115: waveform_sig_loopback =6627;
2116: waveform_sig_loopback =2742;
2117: waveform_sig_loopback =2714;
2118: waveform_sig_loopback =3199;
2119: waveform_sig_loopback =4634;
2120: waveform_sig_loopback =5160;
2121: waveform_sig_loopback =2438;
2122: waveform_sig_loopback =3678;
2123: waveform_sig_loopback =4637;
2124: waveform_sig_loopback =3644;
2125: waveform_sig_loopback =4464;
2126: waveform_sig_loopback =3073;
2127: waveform_sig_loopback =4905;
2128: waveform_sig_loopback =4209;
2129: waveform_sig_loopback =3606;
2130: waveform_sig_loopback =4492;
2131: waveform_sig_loopback =4267;
2132: waveform_sig_loopback =4283;
2133: waveform_sig_loopback =3653;
2134: waveform_sig_loopback =5686;
2135: waveform_sig_loopback =3360;
2136: waveform_sig_loopback =4184;
2137: waveform_sig_loopback =5487;
2138: waveform_sig_loopback =3891;
2139: waveform_sig_loopback =4007;
2140: waveform_sig_loopback =5485;
2141: waveform_sig_loopback =4561;
2142: waveform_sig_loopback =3575;
2143: waveform_sig_loopback =5392;
2144: waveform_sig_loopback =5350;
2145: waveform_sig_loopback =3739;
2146: waveform_sig_loopback =4382;
2147: waveform_sig_loopback =6211;
2148: waveform_sig_loopback =4765;
2149: waveform_sig_loopback =3163;
2150: waveform_sig_loopback =6399;
2151: waveform_sig_loopback =5365;
2152: waveform_sig_loopback =3734;
2153: waveform_sig_loopback =7441;
2154: waveform_sig_loopback =1597;
2155: waveform_sig_loopback =5307;
2156: waveform_sig_loopback =7814;
2157: waveform_sig_loopback =4007;
2158: waveform_sig_loopback =4563;
2159: waveform_sig_loopback =4412;
2160: waveform_sig_loopback =6290;
2161: waveform_sig_loopback =6543;
2162: waveform_sig_loopback =3685;
2163: waveform_sig_loopback =5375;
2164: waveform_sig_loopback =6005;
2165: waveform_sig_loopback =4999;
2166: waveform_sig_loopback =5981;
2167: waveform_sig_loopback =4444;
2168: waveform_sig_loopback =6245;
2169: waveform_sig_loopback =5700;
2170: waveform_sig_loopback =4903;
2171: waveform_sig_loopback =5841;
2172: waveform_sig_loopback =5665;
2173: waveform_sig_loopback =5313;
2174: waveform_sig_loopback =5316;
2175: waveform_sig_loopback =7111;
2176: waveform_sig_loopback =4080;
2177: waveform_sig_loopback =5932;
2178: waveform_sig_loopback =6775;
2179: waveform_sig_loopback =5000;
2180: waveform_sig_loopback =5611;
2181: waveform_sig_loopback =6285;
2182: waveform_sig_loopback =6234;
2183: waveform_sig_loopback =4908;
2184: waveform_sig_loopback =6308;
2185: waveform_sig_loopback =6943;
2186: waveform_sig_loopback =4708;
2187: waveform_sig_loopback =5729;
2188: waveform_sig_loopback =7515;
2189: waveform_sig_loopback =5534;
2190: waveform_sig_loopback =4671;
2191: waveform_sig_loopback =7633;
2192: waveform_sig_loopback =6138;
2193: waveform_sig_loopback =5312;
2194: waveform_sig_loopback =8416;
2195: waveform_sig_loopback =2560;
2196: waveform_sig_loopback =6817;
2197: waveform_sig_loopback =8641;
2198: waveform_sig_loopback =5251;
2199: waveform_sig_loopback =5672;
2200: waveform_sig_loopback =5342;
2201: waveform_sig_loopback =7567;
2202: waveform_sig_loopback =7659;
2203: waveform_sig_loopback =4491;
2204: waveform_sig_loopback =6643;
2205: waveform_sig_loopback =7001;
2206: waveform_sig_loopback =5955;
2207: waveform_sig_loopback =7249;
2208: waveform_sig_loopback =5147;
2209: waveform_sig_loopback =7504;
2210: waveform_sig_loopback =6814;
2211: waveform_sig_loopback =5519;
2212: waveform_sig_loopback =7173;
2213: waveform_sig_loopback =6686;
2214: waveform_sig_loopback =6070;
2215: waveform_sig_loopback =6694;
2216: waveform_sig_loopback =7518;
2217: waveform_sig_loopback =5447;
2218: waveform_sig_loopback =7121;
2219: waveform_sig_loopback =7041;
2220: waveform_sig_loopback =6394;
2221: waveform_sig_loopback =6250;
2222: waveform_sig_loopback =7431;
2223: waveform_sig_loopback =7020;
2224: waveform_sig_loopback =5427;
2225: waveform_sig_loopback =7669;
2226: waveform_sig_loopback =7557;
2227: waveform_sig_loopback =5434;
2228: waveform_sig_loopback =6670;
2229: waveform_sig_loopback =8454;
2230: waveform_sig_loopback =6191;
2231: waveform_sig_loopback =5483;
2232: waveform_sig_loopback =8606;
2233: waveform_sig_loopback =6618;
2234: waveform_sig_loopback =6528;
2235: waveform_sig_loopback =8743;
2236: waveform_sig_loopback =3243;
2237: waveform_sig_loopback =8165;
2238: waveform_sig_loopback =8774;
2239: waveform_sig_loopback =6209;
2240: waveform_sig_loopback =6309;
2241: waveform_sig_loopback =5916;
2242: waveform_sig_loopback =8727;
2243: waveform_sig_loopback =7746;
2244: waveform_sig_loopback =5280;
2245: waveform_sig_loopback =7670;
2246: waveform_sig_loopback =7082;
2247: waveform_sig_loopback =7011;
2248: waveform_sig_loopback =7611;
2249: waveform_sig_loopback =5601;
2250: waveform_sig_loopback =8573;
2251: waveform_sig_loopback =6787;
2252: waveform_sig_loopback =6382;
2253: waveform_sig_loopback =7857;
2254: waveform_sig_loopback =6856;
2255: waveform_sig_loopback =6966;
2256: waveform_sig_loopback =7060;
2257: waveform_sig_loopback =7940;
2258: waveform_sig_loopback =6130;
2259: waveform_sig_loopback =7409;
2260: waveform_sig_loopback =7612;
2261: waveform_sig_loopback =6898;
2262: waveform_sig_loopback =6600;
2263: waveform_sig_loopback =7993;
2264: waveform_sig_loopback =7407;
2265: waveform_sig_loopback =5744;
2266: waveform_sig_loopback =8266;
2267: waveform_sig_loopback =7874;
2268: waveform_sig_loopback =5601;
2269: waveform_sig_loopback =7419;
2270: waveform_sig_loopback =8566;
2271: waveform_sig_loopback =6368;
2272: waveform_sig_loopback =6223;
2273: waveform_sig_loopback =8588;
2274: waveform_sig_loopback =7040;
2275: waveform_sig_loopback =6966;
2276: waveform_sig_loopback =8614;
2277: waveform_sig_loopback =3940;
2278: waveform_sig_loopback =8260;
2279: waveform_sig_loopback =8918;
2280: waveform_sig_loopback =6752;
2281: waveform_sig_loopback =6016;
2282: waveform_sig_loopback =6507;
2283: waveform_sig_loopback =8923;
2284: waveform_sig_loopback =7590;
2285: waveform_sig_loopback =5887;
2286: waveform_sig_loopback =7499;
2287: waveform_sig_loopback =7257;
2288: waveform_sig_loopback =7505;
2289: waveform_sig_loopback =7306;
2290: waveform_sig_loopback =6105;
2291: waveform_sig_loopback =8663;
2292: waveform_sig_loopback =6656;
2293: waveform_sig_loopback =6903;
2294: waveform_sig_loopback =7604;
2295: waveform_sig_loopback =7007;
2296: waveform_sig_loopback =7114;
2297: waveform_sig_loopback =7008;
2298: waveform_sig_loopback =8109;
2299: waveform_sig_loopback =6087;
2300: waveform_sig_loopback =7441;
2301: waveform_sig_loopback =7692;
2302: waveform_sig_loopback =6861;
2303: waveform_sig_loopback =6404;
2304: waveform_sig_loopback =8210;
2305: waveform_sig_loopback =7114;
2306: waveform_sig_loopback =5572;
2307: waveform_sig_loopback =8543;
2308: waveform_sig_loopback =7324;
2309: waveform_sig_loopback =5586;
2310: waveform_sig_loopback =7526;
2311: waveform_sig_loopback =8003;
2312: waveform_sig_loopback =6594;
2313: waveform_sig_loopback =5823;
2314: waveform_sig_loopback =8390;
2315: waveform_sig_loopback =7152;
2316: waveform_sig_loopback =6358;
2317: waveform_sig_loopback =8627;
2318: waveform_sig_loopback =3661;
2319: waveform_sig_loopback =7998;
2320: waveform_sig_loopback =9082;
2321: waveform_sig_loopback =6008;
2322: waveform_sig_loopback =5922;
2323: waveform_sig_loopback =6676;
2324: waveform_sig_loopback =8179;
2325: waveform_sig_loopback =7528;
2326: waveform_sig_loopback =5487;
2327: waveform_sig_loopback =7173;
2328: waveform_sig_loopback =7164;
2329: waveform_sig_loopback =6852;
2330: waveform_sig_loopback =6919;
2331: waveform_sig_loopback =5972;
2332: waveform_sig_loopback =8033;
2333: waveform_sig_loopback =6188;
2334: waveform_sig_loopback =6585;
2335: waveform_sig_loopback =7095;
2336: waveform_sig_loopback =6613;
2337: waveform_sig_loopback =6653;
2338: waveform_sig_loopback =6329;
2339: waveform_sig_loopback =7861;
2340: waveform_sig_loopback =5467;
2341: waveform_sig_loopback =6767;
2342: waveform_sig_loopback =7562;
2343: waveform_sig_loopback =5906;
2344: waveform_sig_loopback =6209;
2345: waveform_sig_loopback =7767;
2346: waveform_sig_loopback =6109;
2347: waveform_sig_loopback =5681;
2348: waveform_sig_loopback =7681;
2349: waveform_sig_loopback =6674;
2350: waveform_sig_loopback =5365;
2351: waveform_sig_loopback =6675;
2352: waveform_sig_loopback =7606;
2353: waveform_sig_loopback =5913;
2354: waveform_sig_loopback =5027;
2355: waveform_sig_loopback =8181;
2356: waveform_sig_loopback =6149;
2357: waveform_sig_loopback =5827;
2358: waveform_sig_loopback =8140;
2359: waveform_sig_loopback =2635;
2360: waveform_sig_loopback =7592;
2361: waveform_sig_loopback =8358;
2362: waveform_sig_loopback =4985;
2363: waveform_sig_loopback =5476;
2364: waveform_sig_loopback =5833;
2365: waveform_sig_loopback =7293;
2366: waveform_sig_loopback =7080;
2367: waveform_sig_loopback =4364;
2368: waveform_sig_loopback =6510;
2369: waveform_sig_loopback =6410;
2370: waveform_sig_loopback =5861;
2371: waveform_sig_loopback =6267;
2372: waveform_sig_loopback =5090;
2373: waveform_sig_loopback =7084;
2374: waveform_sig_loopback =5530;
2375: waveform_sig_loopback =5638;
2376: waveform_sig_loopback =6081;
2377: waveform_sig_loopback =6029;
2378: waveform_sig_loopback =5445;
2379: waveform_sig_loopback =5671;
2380: waveform_sig_loopback =6965;
2381: waveform_sig_loopback =4236;
2382: waveform_sig_loopback =6214;
2383: waveform_sig_loopback =6463;
2384: waveform_sig_loopback =4683;
2385: waveform_sig_loopback =5637;
2386: waveform_sig_loopback =6547;
2387: waveform_sig_loopback =5028;
2388: waveform_sig_loopback =4902;
2389: waveform_sig_loopback =6332;
2390: waveform_sig_loopback =5937;
2391: waveform_sig_loopback =4192;
2392: waveform_sig_loopback =5465;
2393: waveform_sig_loopback =6981;
2394: waveform_sig_loopback =4350;
2395: waveform_sig_loopback =4210;
2396: waveform_sig_loopback =7282;
2397: waveform_sig_loopback =4561;
2398: waveform_sig_loopback =5232;
2399: waveform_sig_loopback =6642;
2400: waveform_sig_loopback =1342;
2401: waveform_sig_loopback =7024;
2402: waveform_sig_loopback =6761;
2403: waveform_sig_loopback =3891;
2404: waveform_sig_loopback =4425;
2405: waveform_sig_loopback =4428;
2406: waveform_sig_loopback =6403;
2407: waveform_sig_loopback =5757;
2408: waveform_sig_loopback =2964;
2409: waveform_sig_loopback =5689;
2410: waveform_sig_loopback =4906;
2411: waveform_sig_loopback =4682;
2412: waveform_sig_loopback =5161;
2413: waveform_sig_loopback =3624;
2414: waveform_sig_loopback =6035;
2415: waveform_sig_loopback =4213;
2416: waveform_sig_loopback =4287;
2417: waveform_sig_loopback =4957;
2418: waveform_sig_loopback =4715;
2419: waveform_sig_loopback =3898;
2420: waveform_sig_loopback =4716;
2421: waveform_sig_loopback =5431;
2422: waveform_sig_loopback =2846;
2423: waveform_sig_loopback =5232;
2424: waveform_sig_loopback =4629;
2425: waveform_sig_loopback =3692;
2426: waveform_sig_loopback =4291;
2427: waveform_sig_loopback =4920;
2428: waveform_sig_loopback =4030;
2429: waveform_sig_loopback =3107;
2430: waveform_sig_loopback =5050;
2431: waveform_sig_loopback =4811;
2432: waveform_sig_loopback =2481;
2433: waveform_sig_loopback =4268;
2434: waveform_sig_loopback =5320;
2435: waveform_sig_loopback =2760;
2436: waveform_sig_loopback =3324;
2437: waveform_sig_loopback =5430;
2438: waveform_sig_loopback =2912;
2439: waveform_sig_loopback =4291;
2440: waveform_sig_loopback =4669;
2441: waveform_sig_loopback =106;
2442: waveform_sig_loopback =5709;
2443: waveform_sig_loopback =4914;
2444: waveform_sig_loopback =2687;
2445: waveform_sig_loopback =2561;
2446: waveform_sig_loopback =3041;
2447: waveform_sig_loopback =5196;
2448: waveform_sig_loopback =3722;
2449: waveform_sig_loopback =1538;
2450: waveform_sig_loopback =4301;
2451: waveform_sig_loopback =3098;
2452: waveform_sig_loopback =3406;
2453: waveform_sig_loopback =3379;
2454: waveform_sig_loopback =1995;
2455: waveform_sig_loopback =4795;
2456: waveform_sig_loopback =2291;
2457: waveform_sig_loopback =2715;
2458: waveform_sig_loopback =3542;
2459: waveform_sig_loopback =2825;
2460: waveform_sig_loopback =2454;
2461: waveform_sig_loopback =3216;
2462: waveform_sig_loopback =3412;
2463: waveform_sig_loopback =1579;
2464: waveform_sig_loopback =3383;
2465: waveform_sig_loopback =2933;
2466: waveform_sig_loopback =2470;
2467: waveform_sig_loopback =2091;
2468: waveform_sig_loopback =3539;
2469: waveform_sig_loopback =2429;
2470: waveform_sig_loopback =1271;
2471: waveform_sig_loopback =3826;
2472: waveform_sig_loopback =2459;
2473: waveform_sig_loopback =867;
2474: waveform_sig_loopback =3172;
2475: waveform_sig_loopback =3106;
2476: waveform_sig_loopback =1314;
2477: waveform_sig_loopback =1470;
2478: waveform_sig_loopback =3755;
2479: waveform_sig_loopback =1435;
2480: waveform_sig_loopback =2333;
2481: waveform_sig_loopback =2937;
2482: waveform_sig_loopback =-1572;
2483: waveform_sig_loopback =4056;
2484: waveform_sig_loopback =3092;
2485: waveform_sig_loopback =935;
2486: waveform_sig_loopback =825;
2487: waveform_sig_loopback =1268;
2488: waveform_sig_loopback =3572;
2489: waveform_sig_loopback =1750;
2490: waveform_sig_loopback =52;
2491: waveform_sig_loopback =2463;
2492: waveform_sig_loopback =1064;
2493: waveform_sig_loopback =2105;
2494: waveform_sig_loopback =1149;
2495: waveform_sig_loopback =455;
2496: waveform_sig_loopback =3056;
2497: waveform_sig_loopback =136;
2498: waveform_sig_loopback =1394;
2499: waveform_sig_loopback =1428;
2500: waveform_sig_loopback =1021;
2501: waveform_sig_loopback =946;
2502: waveform_sig_loopback =1025;
2503: waveform_sig_loopback =1792;
2504: waveform_sig_loopback =-173;
2505: waveform_sig_loopback =1366;
2506: waveform_sig_loopback =1450;
2507: waveform_sig_loopback =131;
2508: waveform_sig_loopback =532;
2509: waveform_sig_loopback =1862;
2510: waveform_sig_loopback =82;
2511: waveform_sig_loopback =-224;
2512: waveform_sig_loopback =1951;
2513: waveform_sig_loopback =523;
2514: waveform_sig_loopback =-886;
2515: waveform_sig_loopback =1190;
2516: waveform_sig_loopback =1331;
2517: waveform_sig_loopback =-583;
2518: waveform_sig_loopback =-454;
2519: waveform_sig_loopback =1920;
2520: waveform_sig_loopback =-480;
2521: waveform_sig_loopback =597;
2522: waveform_sig_loopback =719;
2523: waveform_sig_loopback =-3451;
2524: waveform_sig_loopback =2412;
2525: waveform_sig_loopback =1201;
2526: waveform_sig_loopback =-1120;
2527: waveform_sig_loopback =-1334;
2528: waveform_sig_loopback =-35;
2529: waveform_sig_loopback =1509;
2530: waveform_sig_loopback =-329;
2531: waveform_sig_loopback =-1720;
2532: waveform_sig_loopback =368;
2533: waveform_sig_loopback =-367;
2534: waveform_sig_loopback =-111;
2535: waveform_sig_loopback =-990;
2536: waveform_sig_loopback =-889;
2537: waveform_sig_loopback =708;
2538: waveform_sig_loopback =-1634;
2539: waveform_sig_loopback =-466;
2540: waveform_sig_loopback =-741;
2541: waveform_sig_loopback =-411;
2542: waveform_sig_loopback =-1438;
2543: waveform_sig_loopback =-721;
2544: waveform_sig_loopback =82;
2545: waveform_sig_loopback =-2439;
2546: waveform_sig_loopback =-242;
2547: waveform_sig_loopback =-658;
2548: waveform_sig_loopback =-1776;
2549: waveform_sig_loopback =-1155;
2550: waveform_sig_loopback =-281;
2551: waveform_sig_loopback =-1847;
2552: waveform_sig_loopback =-1944;
2553: waveform_sig_loopback =0;
2554: waveform_sig_loopback =-1553;
2555: waveform_sig_loopback =-2633;
2556: waveform_sig_loopback =-664;
2557: waveform_sig_loopback =-677;
2558: waveform_sig_loopback =-2497;
2559: waveform_sig_loopback =-2357;
2560: waveform_sig_loopback =194;
2561: waveform_sig_loopback =-2539;
2562: waveform_sig_loopback =-1348;
2563: waveform_sig_loopback =-967;
2564: waveform_sig_loopback =-5330;
2565: waveform_sig_loopback =501;
2566: waveform_sig_loopback =-615;
2567: waveform_sig_loopback =-3282;
2568: waveform_sig_loopback =-2723;
2569: waveform_sig_loopback =-2099;
2570: waveform_sig_loopback =-750;
2571: waveform_sig_loopback =-1732;
2572: waveform_sig_loopback =-3873;
2573: waveform_sig_loopback =-1368;
2574: waveform_sig_loopback =-2329;
2575: waveform_sig_loopback =-2181;
2576: waveform_sig_loopback =-2425;
2577: waveform_sig_loopback =-3076;
2578: waveform_sig_loopback =-1222;
2579: waveform_sig_loopback =-3172;
2580: waveform_sig_loopback =-2608;
2581: waveform_sig_loopback =-2420;
2582: waveform_sig_loopback =-2400;
2583: waveform_sig_loopback =-3318;
2584: waveform_sig_loopback =-2260;
2585: waveform_sig_loopback =-2143;
2586: waveform_sig_loopback =-4150;
2587: waveform_sig_loopback =-2011;
2588: waveform_sig_loopback =-2506;
2589: waveform_sig_loopback =-3764;
2590: waveform_sig_loopback =-2850;
2591: waveform_sig_loopback =-2055;
2592: waveform_sig_loopback =-3861;
2593: waveform_sig_loopback =-3450;
2594: waveform_sig_loopback =-2092;
2595: waveform_sig_loopback =-3196;
2596: waveform_sig_loopback =-4355;
2597: waveform_sig_loopback =-2724;
2598: waveform_sig_loopback =-2039;
2599: waveform_sig_loopback =-4600;
2600: waveform_sig_loopback =-3990;
2601: waveform_sig_loopback =-1351;
2602: waveform_sig_loopback =-4853;
2603: waveform_sig_loopback =-2393;
2604: waveform_sig_loopback =-3225;
2605: waveform_sig_loopback =-7181;
2606: waveform_sig_loopback =-590;
2607: waveform_sig_loopback =-2982;
2608: waveform_sig_loopback =-4757;
2609: waveform_sig_loopback =-4423;
2610: waveform_sig_loopback =-4027;
2611: waveform_sig_loopback =-2015;
2612: waveform_sig_loopback =-3842;
2613: waveform_sig_loopback =-5487;
2614: waveform_sig_loopback =-2842;
2615: waveform_sig_loopback =-4297;
2616: waveform_sig_loopback =-3662;
2617: waveform_sig_loopback =-4172;
2618: waveform_sig_loopback =-4719;
2619: waveform_sig_loopback =-2835;
2620: waveform_sig_loopback =-4907;
2621: waveform_sig_loopback =-4267;
2622: waveform_sig_loopback =-3968;
2623: waveform_sig_loopback =-4027;
2624: waveform_sig_loopback =-5156;
2625: waveform_sig_loopback =-3578;
2626: waveform_sig_loopback =-4040;
2627: waveform_sig_loopback =-5734;
2628: waveform_sig_loopback =-3361;
2629: waveform_sig_loopback =-4521;
2630: waveform_sig_loopback =-5052;
2631: waveform_sig_loopback =-4443;
2632: waveform_sig_loopback =-3880;
2633: waveform_sig_loopback =-5146;
2634: waveform_sig_loopback =-5298;
2635: waveform_sig_loopback =-3510;
2636: waveform_sig_loopback =-4731;
2637: waveform_sig_loopback =-6190;
2638: waveform_sig_loopback =-3879;
2639: waveform_sig_loopback =-3800;
2640: waveform_sig_loopback =-6359;
2641: waveform_sig_loopback =-5154;
2642: waveform_sig_loopback =-3088;
2643: waveform_sig_loopback =-6411;
2644: waveform_sig_loopback =-3692;
2645: waveform_sig_loopback =-5211;
2646: waveform_sig_loopback =-8280;
2647: waveform_sig_loopback =-2019;
2648: waveform_sig_loopback =-4868;
2649: waveform_sig_loopback =-5934;
2650: waveform_sig_loopback =-6092;
2651: waveform_sig_loopback =-5398;
2652: waveform_sig_loopback =-3292;
2653: waveform_sig_loopback =-5770;
2654: waveform_sig_loopback =-6663;
2655: waveform_sig_loopback =-4228;
2656: waveform_sig_loopback =-5919;
2657: waveform_sig_loopback =-4800;
2658: waveform_sig_loopback =-5849;
2659: waveform_sig_loopback =-6042;
2660: waveform_sig_loopback =-4105;
2661: waveform_sig_loopback =-6454;
2662: waveform_sig_loopback =-5585;
2663: waveform_sig_loopback =-5252;
2664: waveform_sig_loopback =-5607;
2665: waveform_sig_loopback =-6412;
2666: waveform_sig_loopback =-4746;
2667: waveform_sig_loopback =-5775;
2668: waveform_sig_loopback =-6690;
2669: waveform_sig_loopback =-4841;
2670: waveform_sig_loopback =-5956;
2671: waveform_sig_loopback =-6102;
2672: waveform_sig_loopback =-6164;
2673: waveform_sig_loopback =-4799;
2674: waveform_sig_loopback =-6592;
2675: waveform_sig_loopback =-6718;
2676: waveform_sig_loopback =-4390;
2677: waveform_sig_loopback =-6430;
2678: waveform_sig_loopback =-7260;
2679: waveform_sig_loopback =-4997;
2680: waveform_sig_loopback =-5314;
2681: waveform_sig_loopback =-7435;
2682: waveform_sig_loopback =-6305;
2683: waveform_sig_loopback =-4436;
2684: waveform_sig_loopback =-7595;
2685: waveform_sig_loopback =-4671;
2686: waveform_sig_loopback =-6798;
2687: waveform_sig_loopback =-9165;
2688: waveform_sig_loopback =-3158;
2689: waveform_sig_loopback =-6184;
2690: waveform_sig_loopback =-6904;
2691: waveform_sig_loopback =-7455;
2692: waveform_sig_loopback =-6296;
2693: waveform_sig_loopback =-4304;
2694: waveform_sig_loopback =-7221;
2695: waveform_sig_loopback =-7421;
2696: waveform_sig_loopback =-5429;
2697: waveform_sig_loopback =-7071;
2698: waveform_sig_loopback =-5571;
2699: waveform_sig_loopback =-7318;
2700: waveform_sig_loopback =-6785;
2701: waveform_sig_loopback =-5095;
2702: waveform_sig_loopback =-7819;
2703: waveform_sig_loopback =-6192;
2704: waveform_sig_loopback =-6476;
2705: waveform_sig_loopback =-6561;
2706: waveform_sig_loopback =-7179;
2707: waveform_sig_loopback =-5969;
2708: waveform_sig_loopback =-6561;
2709: waveform_sig_loopback =-7586;
2710: waveform_sig_loopback =-5908;
2711: waveform_sig_loopback =-6694;
2712: waveform_sig_loopback =-7130;
2713: waveform_sig_loopback =-6925;
2714: waveform_sig_loopback =-5643;
2715: waveform_sig_loopback =-7657;
2716: waveform_sig_loopback =-7382;
2717: waveform_sig_loopback =-5216;
2718: waveform_sig_loopback =-7465;
2719: waveform_sig_loopback =-7968;
2720: waveform_sig_loopback =-5691;
2721: waveform_sig_loopback =-6337;
2722: waveform_sig_loopback =-8135;
2723: waveform_sig_loopback =-7035;
2724: waveform_sig_loopback =-5383;
2725: waveform_sig_loopback =-8120;
2726: waveform_sig_loopback =-5573;
2727: waveform_sig_loopback =-7701;
2728: waveform_sig_loopback =-9504;
2729: waveform_sig_loopback =-4197;
2730: waveform_sig_loopback =-6658;
2731: waveform_sig_loopback =-7769;
2732: waveform_sig_loopback =-8284;
2733: waveform_sig_loopback =-6524;
2734: waveform_sig_loopback =-5423;
2735: waveform_sig_loopback =-7726;
2736: waveform_sig_loopback =-7960;
2737: waveform_sig_loopback =-6357;
2738: waveform_sig_loopback =-7404;
2739: waveform_sig_loopback =-6371;
2740: waveform_sig_loopback =-7973;
2741: waveform_sig_loopback =-7091;
2742: waveform_sig_loopback =-6026;
2743: waveform_sig_loopback =-8227;
2744: waveform_sig_loopback =-6677;
2745: waveform_sig_loopback =-7229;
2746: waveform_sig_loopback =-6975;
2747: waveform_sig_loopback =-7752;
2748: waveform_sig_loopback =-6471;
2749: waveform_sig_loopback =-7116;
2750: waveform_sig_loopback =-8078;
2751: waveform_sig_loopback =-6433;
2752: waveform_sig_loopback =-7000;
2753: waveform_sig_loopback =-7830;
2754: waveform_sig_loopback =-7259;
2755: waveform_sig_loopback =-5952;
2756: waveform_sig_loopback =-8466;
2757: waveform_sig_loopback =-7384;
2758: waveform_sig_loopback =-5787;
2759: waveform_sig_loopback =-8033;
2760: waveform_sig_loopback =-7998;
2761: waveform_sig_loopback =-6324;
2762: waveform_sig_loopback =-6603;
2763: waveform_sig_loopback =-8445;
2764: waveform_sig_loopback =-7428;
2765: waveform_sig_loopback =-5508;
2766: waveform_sig_loopback =-8613;
2767: waveform_sig_loopback =-5791;
2768: waveform_sig_loopback =-7995;
2769: waveform_sig_loopback =-9787;
2770: waveform_sig_loopback =-4328;
2771: waveform_sig_loopback =-6879;
2772: waveform_sig_loopback =-8276;
2773: waveform_sig_loopback =-8219;
2774: waveform_sig_loopback =-6731;
2775: waveform_sig_loopback =-5803;
2776: waveform_sig_loopback =-7685;
2777: waveform_sig_loopback =-8318;
2778: waveform_sig_loopback =-6391;
2779: waveform_sig_loopback =-7491;
2780: waveform_sig_loopback =-6730;
2781: waveform_sig_loopback =-7902;
2782: waveform_sig_loopback =-7199;
2783: waveform_sig_loopback =-6271;
2784: waveform_sig_loopback =-8186;
2785: waveform_sig_loopback =-6811;
2786: waveform_sig_loopback =-7319;
2787: waveform_sig_loopback =-6997;
2788: waveform_sig_loopback =-7844;
2789: waveform_sig_loopback =-6453;
2790: waveform_sig_loopback =-7060;
2791: waveform_sig_loopback =-8211;
2792: waveform_sig_loopback =-6265;
2793: waveform_sig_loopback =-6959;
2794: waveform_sig_loopback =-8070;
2795: waveform_sig_loopback =-6761;
2796: waveform_sig_loopback =-6243;
2797: waveform_sig_loopback =-8402;
2798: waveform_sig_loopback =-6979;
2799: waveform_sig_loopback =-6101;
2800: waveform_sig_loopback =-7672;
2801: waveform_sig_loopback =-7948;
2802: waveform_sig_loopback =-6265;
2803: waveform_sig_loopback =-6269;
2804: waveform_sig_loopback =-8601;
2805: waveform_sig_loopback =-7029;
2806: waveform_sig_loopback =-5304;
2807: waveform_sig_loopback =-8677;
2808: waveform_sig_loopback =-5277;
2809: waveform_sig_loopback =-8059;
2810: waveform_sig_loopback =-9503;
2811: waveform_sig_loopback =-3847;
2812: waveform_sig_loopback =-6926;
2813: waveform_sig_loopback =-8024;
2814: waveform_sig_loopback =-7744;
2815: waveform_sig_loopback =-6542;
2816: waveform_sig_loopback =-5414;
2817: waveform_sig_loopback =-7465;
2818: waveform_sig_loopback =-8091;
2819: waveform_sig_loopback =-5817;
2820: waveform_sig_loopback =-7193;
2821: waveform_sig_loopback =-6492;
2822: waveform_sig_loopback =-7381;
2823: waveform_sig_loopback =-6903;
2824: waveform_sig_loopback =-5885;
2825: waveform_sig_loopback =-7676;
2826: waveform_sig_loopback =-6549;
2827: waveform_sig_loopback =-6791;
2828: waveform_sig_loopback =-6498;
2829: waveform_sig_loopback =-7649;
2830: waveform_sig_loopback =-5676;
2831: waveform_sig_loopback =-6845;
2832: waveform_sig_loopback =-7764;
2833: waveform_sig_loopback =-5407;
2834: waveform_sig_loopback =-6953;
2835: waveform_sig_loopback =-7273;
2836: waveform_sig_loopback =-6159;
2837: waveform_sig_loopback =-6032;
2838: waveform_sig_loopback =-7480;
2839: waveform_sig_loopback =-6603;
2840: waveform_sig_loopback =-5457;
2841: waveform_sig_loopback =-7040;
2842: waveform_sig_loopback =-7488;
2843: waveform_sig_loopback =-5368;
2844: waveform_sig_loopback =-5745;
2845: waveform_sig_loopback =-8113;
2846: waveform_sig_loopback =-6053;
2847: waveform_sig_loopback =-4733;
2848: waveform_sig_loopback =-8134;
2849: waveform_sig_loopback =-4246;
2850: waveform_sig_loopback =-7817;
2851: waveform_sig_loopback =-8500;
2852: waveform_sig_loopback =-2905;
2853: waveform_sig_loopback =-6622;
2854: waveform_sig_loopback =-7008;
2855: waveform_sig_loopback =-7001;
2856: waveform_sig_loopback =-5959;
2857: waveform_sig_loopback =-4284;
2858: waveform_sig_loopback =-7029;
2859: waveform_sig_loopback =-7136;
2860: waveform_sig_loopback =-4861;
2861: waveform_sig_loopback =-6756;
2862: waveform_sig_loopback =-5309;
2863: waveform_sig_loopback =-6724;
2864: waveform_sig_loopback =-6055;
2865: waveform_sig_loopback =-4885;
2866: waveform_sig_loopback =-6935;
2867: waveform_sig_loopback =-5644;
2868: waveform_sig_loopback =-5779;
2869: waveform_sig_loopback =-5711;
2870: waveform_sig_loopback =-6686;
2871: waveform_sig_loopback =-4510;
2872: waveform_sig_loopback =-6482;
2873: waveform_sig_loopback =-6444;
2874: waveform_sig_loopback =-4387;
2875: waveform_sig_loopback =-6266;
2876: waveform_sig_loopback =-6125;
2877: waveform_sig_loopback =-5412;
2878: waveform_sig_loopback =-4787;
2879: waveform_sig_loopback =-6372;
2880: waveform_sig_loopback =-6002;
2881: waveform_sig_loopback =-4160;
2882: waveform_sig_loopback =-5974;
2883: waveform_sig_loopback =-6620;
2884: waveform_sig_loopback =-4042;
2885: waveform_sig_loopback =-5031;
2886: waveform_sig_loopback =-6885;
2887: waveform_sig_loopback =-4705;
2888: waveform_sig_loopback =-4221;
2889: waveform_sig_loopback =-6649;
2890: waveform_sig_loopback =-3069;
2891: waveform_sig_loopback =-7146;
2892: waveform_sig_loopback =-6956;
2893: waveform_sig_loopback =-1966;
2894: waveform_sig_loopback =-5450;
2895: waveform_sig_loopback =-5795;
2896: waveform_sig_loopback =-6117;
2897: waveform_sig_loopback =-4528;
2898: waveform_sig_loopback =-3028;
2899: waveform_sig_loopback =-6189;
2900: waveform_sig_loopback =-5710;
2901: waveform_sig_loopback =-3698;
2902: waveform_sig_loopback =-5626;
2903: waveform_sig_loopback =-3819;
2904: waveform_sig_loopback =-5822;
2905: waveform_sig_loopback =-4572;
2906: waveform_sig_loopback =-3511;
2907: waveform_sig_loopback =-6007;
2908: waveform_sig_loopback =-4116;
2909: waveform_sig_loopback =-4425;
2910: waveform_sig_loopback =-4688;
2911: waveform_sig_loopback =-4999;
2912: waveform_sig_loopback =-3432;
2913: waveform_sig_loopback =-5014;
2914: waveform_sig_loopback =-4772;
2915: waveform_sig_loopback =-3594;
2916: waveform_sig_loopback =-4562;
2917: waveform_sig_loopback =-4646;
2918: waveform_sig_loopback =-4165;
2919: waveform_sig_loopback =-3321;
2920: waveform_sig_loopback =-5286;
2921: waveform_sig_loopback =-4288;
2922: waveform_sig_loopback =-2585;
2923: waveform_sig_loopback =-5122;
2924: waveform_sig_loopback =-4898;
2925: waveform_sig_loopback =-2447;
2926: waveform_sig_loopback =-3945;
2927: waveform_sig_loopback =-5255;
2928: waveform_sig_loopback =-3287;
2929: waveform_sig_loopback =-2790;
2930: waveform_sig_loopback =-5003;
2931: waveform_sig_loopback =-1814;
2932: waveform_sig_loopback =-5747;
2933: waveform_sig_loopback =-5065;
2934: waveform_sig_loopback =-719;
2935: waveform_sig_loopback =-3951;
2936: waveform_sig_loopback =-4270;
2937: waveform_sig_loopback =-4658;
2938: waveform_sig_loopback =-2719;
2939: waveform_sig_loopback =-1718;
2940: waveform_sig_loopback =-4734;
2941: waveform_sig_loopback =-3737;
2942: waveform_sig_loopback =-2491;
2943: waveform_sig_loopback =-3955;
2944: waveform_sig_loopback =-2083;
2945: waveform_sig_loopback =-4603;
2946: waveform_sig_loopback =-2578;
2947: waveform_sig_loopback =-2207;
2948: waveform_sig_loopback =-4454;
2949: waveform_sig_loopback =-2117;
2950: waveform_sig_loopback =-3243;
2951: waveform_sig_loopback =-2902;
2952: waveform_sig_loopback =-3191;
2953: waveform_sig_loopback =-2162;
2954: waveform_sig_loopback =-3029;
2955: waveform_sig_loopback =-3344;
2956: waveform_sig_loopback =-1995;
2957: waveform_sig_loopback =-2574;
2958: waveform_sig_loopback =-3470;
2959: waveform_sig_loopback =-2044;
2960: waveform_sig_loopback =-1809;
2961: waveform_sig_loopback =-3794;
2962: waveform_sig_loopback =-2235;
2963: waveform_sig_loopback =-1192;
2964: waveform_sig_loopback =-3362;
2965: waveform_sig_loopback =-3097;
2966: waveform_sig_loopback =-768;
2967: waveform_sig_loopback =-2287;
2968: waveform_sig_loopback =-3480;
2969: waveform_sig_loopback =-1523;
2970: waveform_sig_loopback =-1188;
2971: waveform_sig_loopback =-3076;
2972: waveform_sig_loopback =-259;
2973: waveform_sig_loopback =-4005;
2974: waveform_sig_loopback =-3087;
2975: waveform_sig_loopback =826;
2976: waveform_sig_loopback =-1925;
2977: waveform_sig_loopback =-2784;
2978: waveform_sig_loopback =-2825;
2979: waveform_sig_loopback =-579;
2980: waveform_sig_loopback =-438;
2981: waveform_sig_loopback =-2679;
2982: waveform_sig_loopback =-1936;
2983: waveform_sig_loopback =-1024;
2984: waveform_sig_loopback =-1650;
2985: waveform_sig_loopback =-805;
2986: waveform_sig_loopback =-2610;
2987: waveform_sig_loopback =-482;
2988: waveform_sig_loopback =-979;
2989: waveform_sig_loopback =-2052;
2990: waveform_sig_loopback =-619;
2991: waveform_sig_loopback =-1487;
2992: waveform_sig_loopback =-736;
2993: waveform_sig_loopback =-1840;
2994: waveform_sig_loopback =86;
2995: waveform_sig_loopback =-1431;
2996: waveform_sig_loopback =-1571;
2997: waveform_sig_loopback =132;
2998: waveform_sig_loopback =-1044;
2999: waveform_sig_loopback =-1442;
3000: waveform_sig_loopback =-227;
3001: waveform_sig_loopback =-24;
3002: waveform_sig_loopback =-1977;
3003: waveform_sig_loopback =-248;
3004: waveform_sig_loopback =623;
3005: waveform_sig_loopback =-1723;
3006: waveform_sig_loopback =-869;
3007: waveform_sig_loopback =786;
3008: waveform_sig_loopback =-369;
3009: waveform_sig_loopback =-1493;
3010: waveform_sig_loopback =63;
3011: waveform_sig_loopback =1082;
3012: waveform_sig_loopback =-1545;
3013: waveform_sig_loopback =1681;
3014: waveform_sig_loopback =-2057;
3015: waveform_sig_loopback =-1504;
3016: waveform_sig_loopback =3147;
3017: waveform_sig_loopback =-356;
3018: waveform_sig_loopback =-1137;
3019: waveform_sig_loopback =-361;
3020: waveform_sig_loopback =796;
3021: waveform_sig_loopback =1645;
3022: waveform_sig_loopback =-745;
3023: waveform_sig_loopback =-372;
3024: waveform_sig_loopback =1253;
3025: waveform_sig_loopback =10;
3026: waveform_sig_loopback =1027;
3027: waveform_sig_loopback =-448;
3028: waveform_sig_loopback =1117;
3029: waveform_sig_loopback =1002;
3030: waveform_sig_loopback =-104;
3031: waveform_sig_loopback =1052;
3032: waveform_sig_loopback =708;
3033: waveform_sig_loopback =899;
3034: waveform_sig_loopback =87;
3035: waveform_sig_loopback =2092;
3036: waveform_sig_loopback =234;
3037: waveform_sig_loopback =420;
3038: waveform_sig_loopback =2041;
3039: waveform_sig_loopback =776;
3040: waveform_sig_loopback =362;
3041: waveform_sig_loopback =1920;
3042: waveform_sig_loopback =1568;
3043: waveform_sig_loopback =19;
3044: waveform_sig_loopback =1837;
3045: waveform_sig_loopback =2171;
3046: waveform_sig_loopback =479;
3047: waveform_sig_loopback =878;
3048: waveform_sig_loopback =2680;
3049: waveform_sig_loopback =1785;
3050: waveform_sig_loopback =-97;
3051: waveform_sig_loopback =2433;
3052: waveform_sig_loopback =2799;
3053: waveform_sig_loopback =68;
3054: waveform_sig_loopback =4147;
3055: waveform_sig_loopback =-906;
3056: waveform_sig_loopback =874;
3057: waveform_sig_loopback =5188;
3058: waveform_sig_loopback =861;
3059: waveform_sig_loopback =1262;
3060: waveform_sig_loopback =1305;
3061: waveform_sig_loopback =2649;
3062: waveform_sig_loopback =3805;
3063: waveform_sig_loopback =580;
3064: waveform_sig_loopback =1911;
3065: waveform_sig_loopback =3081;
3066: waveform_sig_loopback =1656;
3067: waveform_sig_loopback =3089;
3068: waveform_sig_loopback =1234;
3069: waveform_sig_loopback =3062;
3070: waveform_sig_loopback =2837;
3071: waveform_sig_loopback =1681;
3072: waveform_sig_loopback =2931;
3073: waveform_sig_loopback =2623;
3074: waveform_sig_loopback =2628;
3075: waveform_sig_loopback =1853;
3076: waveform_sig_loopback =4148;
3077: waveform_sig_loopback =1744;
3078: waveform_sig_loopback =2421;
3079: waveform_sig_loopback =3984;
3080: waveform_sig_loopback =2137;
3081: waveform_sig_loopback =2638;
3082: waveform_sig_loopback =3523;
3083: waveform_sig_loopback =3200;
3084: waveform_sig_loopback =2185;
3085: waveform_sig_loopback =3217;
3086: waveform_sig_loopback =4269;
3087: waveform_sig_loopback =2124;
3088: waveform_sig_loopback =2474;
3089: waveform_sig_loopback =4922;
3090: waveform_sig_loopback =3003;
3091: waveform_sig_loopback =1810;
3092: waveform_sig_loopback =4565;
3093: waveform_sig_loopback =3952;
3094: waveform_sig_loopback =2297;
3095: waveform_sig_loopback =5727;
3096: waveform_sig_loopback =540;
3097: waveform_sig_loopback =3236;
3098: waveform_sig_loopback =6412;
3099: waveform_sig_loopback =2802;
3100: waveform_sig_loopback =3034;
3101: waveform_sig_loopback =2741;
3102: waveform_sig_loopback =4745;
3103: waveform_sig_loopback =5300;
3104: waveform_sig_loopback =2236;
3105: waveform_sig_loopback =3790;
3106: waveform_sig_loopback =4618;
3107: waveform_sig_loopback =3451;
3108: waveform_sig_loopback =4826;
3109: waveform_sig_loopback =2755;
3110: waveform_sig_loopback =4862;
3111: waveform_sig_loopback =4577;
3112: waveform_sig_loopback =3208;
3113: waveform_sig_loopback =4661;
3114: waveform_sig_loopback =4363;
3115: waveform_sig_loopback =4009;
3116: waveform_sig_loopback =3905;
3117: waveform_sig_loopback =5580;
3118: waveform_sig_loopback =3211;
3119: waveform_sig_loopback =4546;
3120: waveform_sig_loopback =5072;
3121: waveform_sig_loopback =4099;
3122: waveform_sig_loopback =4161;
3123: waveform_sig_loopback =4935;
3124: waveform_sig_loopback =5232;
3125: waveform_sig_loopback =3221;
3126: waveform_sig_loopback =5115;
3127: waveform_sig_loopback =5879;
3128: waveform_sig_loopback =3365;
3129: waveform_sig_loopback =4418;
3130: waveform_sig_loopback =6315;
3131: waveform_sig_loopback =4478;
3132: waveform_sig_loopback =3521;
3133: waveform_sig_loopback =6098;
3134: waveform_sig_loopback =5277;
3135: waveform_sig_loopback =4040;
3136: waveform_sig_loopback =7104;
3137: waveform_sig_loopback =1889;
3138: waveform_sig_loopback =5133;
3139: waveform_sig_loopback =7612;
3140: waveform_sig_loopback =4398;
3141: waveform_sig_loopback =4471;
3142: waveform_sig_loopback =4146;
3143: waveform_sig_loopback =6524;
3144: waveform_sig_loopback =6469;
3145: waveform_sig_loopback =3620;
3146: waveform_sig_loopback =5519;
3147: waveform_sig_loopback =5732;
3148: waveform_sig_loopback =5072;
3149: waveform_sig_loopback =6195;
3150: waveform_sig_loopback =3979;
3151: waveform_sig_loopback =6627;
3152: waveform_sig_loopback =5664;
3153: waveform_sig_loopback =4600;
3154: waveform_sig_loopback =6256;
3155: waveform_sig_loopback =5418;
3156: waveform_sig_loopback =5447;
3157: waveform_sig_loopback =5378;
3158: waveform_sig_loopback =6651;
3159: waveform_sig_loopback =4780;
3160: waveform_sig_loopback =5801;
3161: waveform_sig_loopback =6269;
3162: waveform_sig_loopback =5629;
3163: waveform_sig_loopback =5152;
3164: waveform_sig_loopback =6450;
3165: waveform_sig_loopback =6488;
3166: waveform_sig_loopback =4322;
3167: waveform_sig_loopback =6753;
3168: waveform_sig_loopback =6829;
3169: waveform_sig_loopback =4630;
3170: waveform_sig_loopback =5935;
3171: waveform_sig_loopback =7297;
3172: waveform_sig_loopback =5700;
3173: waveform_sig_loopback =4822;
3174: waveform_sig_loopback =7287;
3175: waveform_sig_loopback =6471;
3176: waveform_sig_loopback =5372;
3177: waveform_sig_loopback =8056;
3178: waveform_sig_loopback =3100;
3179: waveform_sig_loopback =6465;
3180: waveform_sig_loopback =8562;
3181: waveform_sig_loopback =5715;
3182: waveform_sig_loopback =5360;
3183: waveform_sig_loopback =5400;
3184: waveform_sig_loopback =7774;
3185: waveform_sig_loopback =7249;
3186: waveform_sig_loopback =4973;
3187: waveform_sig_loopback =6538;
3188: waveform_sig_loopback =6648;
3189: waveform_sig_loopback =6505;
3190: waveform_sig_loopback =6877;
3191: waveform_sig_loopback =5191;
3192: waveform_sig_loopback =7810;
3193: waveform_sig_loopback =6311;
3194: waveform_sig_loopback =5966;
3195: waveform_sig_loopback =7046;
3196: waveform_sig_loopback =6462;
3197: waveform_sig_loopback =6629;
3198: waveform_sig_loopback =6134;
3199: waveform_sig_loopback =7786;
3200: waveform_sig_loopback =5661;
3201: waveform_sig_loopback =6657;
3202: waveform_sig_loopback =7365;
3203: waveform_sig_loopback =6491;
3204: waveform_sig_loopback =6036;
3205: waveform_sig_loopback =7554;
3206: waveform_sig_loopback =7173;
3207: waveform_sig_loopback =5208;
3208: waveform_sig_loopback =7924;
3209: waveform_sig_loopback =7415;
3210: waveform_sig_loopback =5486;
3211: waveform_sig_loopback =6987;
3212: waveform_sig_loopback =7878;
3213: waveform_sig_loopback =6752;
3214: waveform_sig_loopback =5466;
3215: waveform_sig_loopback =8103;
3216: waveform_sig_loopback =7390;
3217: waveform_sig_loopback =5930;
3218: waveform_sig_loopback =8971;
3219: waveform_sig_loopback =3700;
3220: waveform_sig_loopback =7290;
3221: waveform_sig_loopback =9485;
3222: waveform_sig_loopback =6039;
3223: waveform_sig_loopback =5885;
3224: waveform_sig_loopback =6594;
3225: waveform_sig_loopback =8260;
3226: waveform_sig_loopback =7766;
3227: waveform_sig_loopback =5512;
3228: waveform_sig_loopback =7269;
3229: waveform_sig_loopback =7527;
3230: waveform_sig_loopback =6880;
3231: waveform_sig_loopback =7221;
3232: waveform_sig_loopback =6225;
3233: waveform_sig_loopback =8299;
3234: waveform_sig_loopback =6696;
3235: waveform_sig_loopback =6676;
3236: waveform_sig_loopback =7451;
3237: waveform_sig_loopback =7205;
3238: waveform_sig_loopback =7008;
3239: waveform_sig_loopback =6500;
3240: waveform_sig_loopback =8580;
3241: waveform_sig_loopback =5978;
3242: waveform_sig_loopback =7075;
3243: waveform_sig_loopback =8050;
3244: waveform_sig_loopback =6667;
3245: waveform_sig_loopback =6641;
3246: waveform_sig_loopback =8043;
3247: waveform_sig_loopback =7179;
3248: waveform_sig_loopback =6075;
3249: waveform_sig_loopback =8135;
3250: waveform_sig_loopback =7620;
3251: waveform_sig_loopback =6093;
3252: waveform_sig_loopback =7195;
3253: waveform_sig_loopback =8389;
3254: waveform_sig_loopback =6923;
3255: waveform_sig_loopback =5689;
3256: waveform_sig_loopback =8758;
3257: waveform_sig_loopback =7395;
3258: waveform_sig_loopback =6243;
3259: waveform_sig_loopback =9354;
3260: waveform_sig_loopback =3736;
3261: waveform_sig_loopback =7829;
3262: waveform_sig_loopback =9645;
3263: waveform_sig_loopback =6207;
3264: waveform_sig_loopback =6372;
3265: waveform_sig_loopback =6704;
3266: waveform_sig_loopback =8249;
3267: waveform_sig_loopback =8284;
3268: waveform_sig_loopback =5708;
3269: waveform_sig_loopback =7229;
3270: waveform_sig_loopback =7802;
3271: waveform_sig_loopback =6914;
3272: waveform_sig_loopback =7596;
3273: waveform_sig_loopback =6249;
3274: waveform_sig_loopback =8101;
3275: waveform_sig_loopback =7197;
3276: waveform_sig_loopback =6668;
3277: waveform_sig_loopback =7401;
3278: waveform_sig_loopback =7427;
3279: waveform_sig_loopback =6852;
3280: waveform_sig_loopback =6852;
3281: waveform_sig_loopback =8455;
3282: waveform_sig_loopback =5786;
3283: waveform_sig_loopback =7437;
3284: waveform_sig_loopback =7900;
3285: waveform_sig_loopback =6461;
3286: waveform_sig_loopback =6809;
3287: waveform_sig_loopback =8001;
3288: waveform_sig_loopback =6996;
3289: waveform_sig_loopback =6143;
3290: waveform_sig_loopback =7912;
3291: waveform_sig_loopback =7648;
3292: waveform_sig_loopback =5971;
3293: waveform_sig_loopback =6912;
3294: waveform_sig_loopback =8536;
3295: waveform_sig_loopback =6555;
3296: waveform_sig_loopback =5575;
3297: waveform_sig_loopback =8808;
3298: waveform_sig_loopback =6842;
3299: waveform_sig_loopback =6432;
3300: waveform_sig_loopback =9048;
3301: waveform_sig_loopback =3189;
3302: waveform_sig_loopback =8123;
3303: waveform_sig_loopback =9174;
3304: waveform_sig_loopback =5801;
3305: waveform_sig_loopback =6320;
3306: waveform_sig_loopback =6253;
3307: waveform_sig_loopback =8182;
3308: waveform_sig_loopback =7979;
3309: waveform_sig_loopback =5059;
3310: waveform_sig_loopback =7310;
3311: waveform_sig_loopback =7256;
3312: waveform_sig_loopback =6504;
3313: waveform_sig_loopback =7454;
3314: waveform_sig_loopback =5622;
3315: waveform_sig_loopback =7899;
3316: waveform_sig_loopback =6791;
3317: waveform_sig_loopback =6050;
3318: waveform_sig_loopback =7241;
3319: waveform_sig_loopback =6906;
3320: waveform_sig_loopback =6265;
3321: waveform_sig_loopback =6682;
3322: waveform_sig_loopback =7758;
3323: waveform_sig_loopback =5329;
3324: waveform_sig_loopback =7129;
3325: waveform_sig_loopback =7183;
3326: waveform_sig_loopback =6046;
3327: waveform_sig_loopback =6352;
3328: waveform_sig_loopback =7331;
3329: waveform_sig_loopback =6524;
3330: waveform_sig_loopback =5521;
3331: waveform_sig_loopback =7257;
3332: waveform_sig_loopback =7234;
3333: waveform_sig_loopback =5151;
3334: waveform_sig_loopback =6367;
3335: waveform_sig_loopback =8092;
3336: waveform_sig_loopback =5481;
3337: waveform_sig_loopback =5285;
3338: waveform_sig_loopback =8149;
3339: waveform_sig_loopback =5794;
3340: waveform_sig_loopback =6281;
3341: waveform_sig_loopback =7836;
3342: waveform_sig_loopback =2584;
3343: waveform_sig_loopback =7836;
3344: waveform_sig_loopback =7960;
3345: waveform_sig_loopback =5358;
3346: waveform_sig_loopback =5440;
3347: waveform_sig_loopback =5428;
3348: waveform_sig_loopback =7771;
3349: waveform_sig_loopback =6848;
3350: waveform_sig_loopback =4307;
3351: waveform_sig_loopback =6743;
3352: waveform_sig_loopback =6130;
3353: waveform_sig_loopback =5931;
3354: waveform_sig_loopback =6452;
3355: waveform_sig_loopback =4689;
3356: waveform_sig_loopback =7319;
3357: waveform_sig_loopback =5646;
3358: waveform_sig_loopback =5304;
3359: waveform_sig_loopback =6373;
3360: waveform_sig_loopback =5895;
3361: waveform_sig_loopback =5313;
3362: waveform_sig_loopback =5993;
3363: waveform_sig_loopback =6595;
3364: waveform_sig_loopback =4428;
3365: waveform_sig_loopback =6423;
3366: waveform_sig_loopback =5909;
3367: waveform_sig_loopback =5377;
3368: waveform_sig_loopback =5246;
3369: waveform_sig_loopback =6329;
3370: waveform_sig_loopback =5753;
3371: waveform_sig_loopback =4197;
3372: waveform_sig_loopback =6647;
3373: waveform_sig_loopback =6066;
3374: waveform_sig_loopback =3885;
3375: waveform_sig_loopback =5840;
3376: waveform_sig_loopback =6679;
3377: waveform_sig_loopback =4474;
3378: waveform_sig_loopback =4425;
3379: waveform_sig_loopback =6873;
3380: waveform_sig_loopback =4849;
3381: waveform_sig_loopback =5207;
3382: waveform_sig_loopback =6582;
3383: waveform_sig_loopback =1549;
3384: waveform_sig_loopback =6761;
3385: waveform_sig_loopback =6752;
3386: waveform_sig_loopback =4233;
3387: waveform_sig_loopback =4173;
3388: waveform_sig_loopback =4318;
3389: waveform_sig_loopback =6701;
3390: waveform_sig_loopback =5445;
3391: waveform_sig_loopback =3154;
3392: waveform_sig_loopback =5687;
3393: waveform_sig_loopback =4627;
3394: waveform_sig_loopback =5009;
3395: waveform_sig_loopback =5049;
3396: waveform_sig_loopback =3419;
3397: waveform_sig_loopback =6364;
3398: waveform_sig_loopback =3950;
3399: waveform_sig_loopback =4287;
3400: waveform_sig_loopback =5170;
3401: waveform_sig_loopback =4275;
3402: waveform_sig_loopback =4389;
3403: waveform_sig_loopback =4471;
3404: waveform_sig_loopback =5200;
3405: waveform_sig_loopback =3395;
3406: waveform_sig_loopback =4709;
3407: waveform_sig_loopback =4891;
3408: waveform_sig_loopback =3851;
3409: waveform_sig_loopback =3785;
3410: waveform_sig_loopback =5257;
3411: waveform_sig_loopback =4070;
3412: waveform_sig_loopback =2900;
3413: waveform_sig_loopback =5357;
3414: waveform_sig_loopback =4446;
3415: waveform_sig_loopback =2475;
3416: waveform_sig_loopback =4600;
3417: waveform_sig_loopback =4984;
3418: waveform_sig_loopback =3155;
3419: waveform_sig_loopback =3043;
3420: waveform_sig_loopback =5300;
3421: waveform_sig_loopback =3465;
3422: waveform_sig_loopback =3769;
3423: waveform_sig_loopback =4931;
3424: waveform_sig_loopback =196;
3425: waveform_sig_loopback =5336;
3426: waveform_sig_loopback =5158;
3427: waveform_sig_loopback =2784;
3428: waveform_sig_loopback =2443;
3429: waveform_sig_loopback =3070;
3430: waveform_sig_loopback =5195;
3431: waveform_sig_loopback =3570;
3432: waveform_sig_loopback =1987;
3433: waveform_sig_loopback =3909;
3434: waveform_sig_loopback =3105;
3435: waveform_sig_loopback =3712;
3436: waveform_sig_loopback =2954;
3437: waveform_sig_loopback =2328;
3438: waveform_sig_loopback =4612;
3439: waveform_sig_loopback =2136;
3440: waveform_sig_loopback =3145;
3441: waveform_sig_loopback =3121;
3442: waveform_sig_loopback =2979;
3443: waveform_sig_loopback =2733;
3444: waveform_sig_loopback =2650;
3445: waveform_sig_loopback =3889;
3446: waveform_sig_loopback =1482;
3447: waveform_sig_loopback =3181;
3448: waveform_sig_loopback =3315;
3449: waveform_sig_loopback =2011;
3450: waveform_sig_loopback =2343;
3451: waveform_sig_loopback =3550;
3452: waveform_sig_loopback =2177;
3453: waveform_sig_loopback =1464;
3454: waveform_sig_loopback =3673;
3455: waveform_sig_loopback =2570;
3456: waveform_sig_loopback =901;
3457: waveform_sig_loopback =2949;
3458: waveform_sig_loopback =3167;
3459: waveform_sig_loopback =1413;
3460: waveform_sig_loopback =1302;
3461: waveform_sig_loopback =3545;
3462: waveform_sig_loopback =1824;
3463: waveform_sig_loopback =1882;
3464: waveform_sig_loopback =3186;
3465: waveform_sig_loopback =-1437;
3466: waveform_sig_loopback =3402;
3467: waveform_sig_loopback =3774;
3468: waveform_sig_loopback =645;
3469: waveform_sig_loopback =696;
3470: waveform_sig_loopback =1714;
3471: waveform_sig_loopback =2853;
3472: waveform_sig_loopback =2290;
3473: waveform_sig_loopback =-4;
3474: waveform_sig_loopback =2057;
3475: waveform_sig_loopback =1666;
3476: waveform_sig_loopback =1495;
3477: waveform_sig_loopback =1461;
3478: waveform_sig_loopback =617;
3479: waveform_sig_loopback =2510;
3480: waveform_sig_loopback =676;
3481: waveform_sig_loopback =1131;
3482: waveform_sig_loopback =1325;
3483: waveform_sig_loopback =1290;
3484: waveform_sig_loopback =685;
3485: waveform_sig_loopback =1107;
3486: waveform_sig_loopback =1888;
3487: waveform_sig_loopback =-339;
3488: waveform_sig_loopback =1403;
3489: waveform_sig_loopback =1491;
3490: waveform_sig_loopback =69;
3491: waveform_sig_loopback =515;
3492: waveform_sig_loopback =1912;
3493: waveform_sig_loopback =-63;
3494: waveform_sig_loopback =12;
3495: waveform_sig_loopback =1674;
3496: waveform_sig_loopback =517;
3497: waveform_sig_loopback =-563;
3498: waveform_sig_loopback =702;
3499: waveform_sig_loopback =1644;
3500: waveform_sig_loopback =-539;
3501: waveform_sig_loopback =-758;
3502: waveform_sig_loopback =2222;
3503: waveform_sig_loopback =-611;
3504: waveform_sig_loopback =325;
3505: waveform_sig_loopback =1353;
3506: waveform_sig_loopback =-3743;
3507: waveform_sig_loopback =2186;
3508: waveform_sig_loopback =1502;
3509: waveform_sig_loopback =-1450;
3510: waveform_sig_loopback =-701;
3511: waveform_sig_loopback =-506;
3512: waveform_sig_loopback =1159;
3513: waveform_sig_loopback =418;
3514: waveform_sig_loopback =-2121;
3515: waveform_sig_loopback =608;
3516: waveform_sig_loopback =-493;
3517: waveform_sig_loopback =-434;
3518: waveform_sig_loopback =-241;
3519: waveform_sig_loopback =-1412;
3520: waveform_sig_loopback =675;
3521: waveform_sig_loopback =-1253;
3522: waveform_sig_loopback =-829;
3523: waveform_sig_loopback =-417;
3524: waveform_sig_loopback =-612;
3525: waveform_sig_loopback =-1338;
3526: waveform_sig_loopback =-673;
3527: waveform_sig_loopback =30;
3528: waveform_sig_loopback =-2426;
3529: waveform_sig_loopback =-188;
3530: waveform_sig_loopback =-504;
3531: waveform_sig_loopback =-2037;
3532: waveform_sig_loopback =-871;
3533: waveform_sig_loopback =-470;
3534: waveform_sig_loopback =-1687;
3535: waveform_sig_loopback =-1718;
3536: waveform_sig_loopback =-545;
3537: waveform_sig_loopback =-930;
3538: waveform_sig_loopback =-2834;
3539: waveform_sig_loopback =-945;
3540: waveform_sig_loopback =-57;
3541: waveform_sig_loopback =-2858;
3542: waveform_sig_loopback =-2131;
3543: waveform_sig_loopback =287;
3544: waveform_sig_loopback =-2809;
3545: waveform_sig_loopback =-931;
3546: waveform_sig_loopback =-1042;
3547: waveform_sig_loopback =-5453;
3548: waveform_sig_loopback =758;
3549: waveform_sig_loopback =-875;
3550: waveform_sig_loopback =-2926;
3551: waveform_sig_loopback =-2709;
3552: waveform_sig_loopback =-2494;
3553: waveform_sig_loopback =-256;
3554: waveform_sig_loopback =-1894;
3555: waveform_sig_loopback =-3916;
3556: waveform_sig_loopback =-1114;
3557: waveform_sig_loopback =-2531;
3558: waveform_sig_loopback =-2009;
3559: waveform_sig_loopback =-2314;
3560: waveform_sig_loopback =-3347;
3561: waveform_sig_loopback =-981;
3562: waveform_sig_loopback =-3160;
3563: waveform_sig_loopback =-2695;
3564: waveform_sig_loopback =-2256;
3565: waveform_sig_loopback =-2407;
3566: waveform_sig_loopback =-3362;
3567: waveform_sig_loopback =-2147;
3568: waveform_sig_loopback =-2187;
3569: waveform_sig_loopback =-4189;
3570: waveform_sig_loopback =-1649;
3571: waveform_sig_loopback =-3148;
3572: waveform_sig_loopback =-3230;
3573: waveform_sig_loopback =-2877;
3574: waveform_sig_loopback =-2400;
3575: waveform_sig_loopback =-3360;
3576: waveform_sig_loopback =-4158;
3577: waveform_sig_loopback =-1555;
3578: waveform_sig_loopback =-3087;
3579: waveform_sig_loopback =-4893;
3580: waveform_sig_loopback =-2322;
3581: waveform_sig_loopback =-2171;
3582: waveform_sig_loopback =-4591;
3583: waveform_sig_loopback =-3905;
3584: waveform_sig_loopback =-1676;
3585: waveform_sig_loopback =-4516;
3586: waveform_sig_loopback =-2578;
3587: waveform_sig_loopback =-3307;
3588: waveform_sig_loopback =-7013;
3589: waveform_sig_loopback =-811;
3590: waveform_sig_loopback =-3004;
3591: waveform_sig_loopback =-4537;
3592: waveform_sig_loopback =-4598;
3593: waveform_sig_loopback =-4061;
3594: waveform_sig_loopback =-1845;
3595: waveform_sig_loopback =-4067;
3596: waveform_sig_loopback =-5379;
3597: waveform_sig_loopback =-2709;
3598: waveform_sig_loopback =-4590;
3599: waveform_sig_loopback =-3390;
3600: waveform_sig_loopback =-4264;
3601: waveform_sig_loopback =-4895;
3602: waveform_sig_loopback =-2475;
3603: waveform_sig_loopback =-5244;
3604: waveform_sig_loopback =-4100;
3605: waveform_sig_loopback =-3890;
3606: waveform_sig_loopback =-4358;
3607: waveform_sig_loopback =-4692;
3608: waveform_sig_loopback =-3780;
3609: waveform_sig_loopback =-4116;
3610: waveform_sig_loopback =-5474;
3611: waveform_sig_loopback =-3598;
3612: waveform_sig_loopback =-4366;
3613: waveform_sig_loopback =-4873;
3614: waveform_sig_loopback =-4918;
3615: waveform_sig_loopback =-3530;
3616: waveform_sig_loopback =-5034;
3617: waveform_sig_loopback =-5668;
3618: waveform_sig_loopback =-3125;
3619: waveform_sig_loopback =-5040;
3620: waveform_sig_loopback =-6115;
3621: waveform_sig_loopback =-3677;
3622: waveform_sig_loopback =-4162;
3623: waveform_sig_loopback =-5961;
3624: waveform_sig_loopback =-5297;
3625: waveform_sig_loopback =-3293;
3626: waveform_sig_loopback =-5961;
3627: waveform_sig_loopback =-4090;
3628: waveform_sig_loopback =-4896;
3629: waveform_sig_loopback =-8258;
3630: waveform_sig_loopback =-2489;
3631: waveform_sig_loopback =-4386;
3632: waveform_sig_loopback =-5971;
3633: waveform_sig_loopback =-6380;
3634: waveform_sig_loopback =-5214;
3635: waveform_sig_loopback =-3460;
3636: waveform_sig_loopback =-5659;
3637: waveform_sig_loopback =-6545;
3638: waveform_sig_loopback =-4497;
3639: waveform_sig_loopback =-5815;
3640: waveform_sig_loopback =-4696;
3641: waveform_sig_loopback =-6011;
3642: waveform_sig_loopback =-5941;
3643: waveform_sig_loopback =-4049;
3644: waveform_sig_loopback =-6662;
3645: waveform_sig_loopback =-5249;
3646: waveform_sig_loopback =-5495;
3647: waveform_sig_loopback =-5602;
3648: waveform_sig_loopback =-6064;
3649: waveform_sig_loopback =-5299;
3650: waveform_sig_loopback =-5308;
3651: waveform_sig_loopback =-6765;
3652: waveform_sig_loopback =-5169;
3653: waveform_sig_loopback =-5429;
3654: waveform_sig_loopback =-6471;
3655: waveform_sig_loopback =-6100;
3656: waveform_sig_loopback =-4595;
3657: waveform_sig_loopback =-6885;
3658: waveform_sig_loopback =-6516;
3659: waveform_sig_loopback =-4487;
3660: waveform_sig_loopback =-6472;
3661: waveform_sig_loopback =-7081;
3662: waveform_sig_loopback =-5196;
3663: waveform_sig_loopback =-5304;
3664: waveform_sig_loopback =-7175;
3665: waveform_sig_loopback =-6639;
3666: waveform_sig_loopback =-4353;
3667: waveform_sig_loopback =-7298;
3668: waveform_sig_loopback =-5220;
3669: waveform_sig_loopback =-6224;
3670: waveform_sig_loopback =-9357;
3671: waveform_sig_loopback =-3554;
3672: waveform_sig_loopback =-5598;
3673: waveform_sig_loopback =-7275;
3674: waveform_sig_loopback =-7350;
3675: waveform_sig_loopback =-6135;
3676: waveform_sig_loopback =-4789;
3677: waveform_sig_loopback =-6677;
3678: waveform_sig_loopback =-7582;
3679: waveform_sig_loopback =-5661;
3680: waveform_sig_loopback =-6678;
3681: waveform_sig_loopback =-5943;
3682: waveform_sig_loopback =-7094;
3683: waveform_sig_loopback =-6688;
3684: waveform_sig_loopback =-5427;
3685: waveform_sig_loopback =-7528;
3686: waveform_sig_loopback =-6238;
3687: waveform_sig_loopback =-6645;
3688: waveform_sig_loopback =-6319;
3689: waveform_sig_loopback =-7264;
3690: waveform_sig_loopback =-6151;
3691: waveform_sig_loopback =-6181;
3692: waveform_sig_loopback =-7963;
3693: waveform_sig_loopback =-5845;
3694: waveform_sig_loopback =-6393;
3695: waveform_sig_loopback =-7586;
3696: waveform_sig_loopback =-6611;
3697: waveform_sig_loopback =-5779;
3698: waveform_sig_loopback =-7762;
3699: waveform_sig_loopback =-7095;
3700: waveform_sig_loopback =-5643;
3701: waveform_sig_loopback =-7155;
3702: waveform_sig_loopback =-7921;
3703: waveform_sig_loopback =-6067;
3704: waveform_sig_loopback =-5956;
3705: waveform_sig_loopback =-8188;
3706: waveform_sig_loopback =-7276;
3707: waveform_sig_loopback =-5078;
3708: waveform_sig_loopback =-8299;
3709: waveform_sig_loopback =-5719;
3710: waveform_sig_loopback =-7213;
3711: waveform_sig_loopback =-10016;
3712: waveform_sig_loopback =-4088;
3713: waveform_sig_loopback =-6460;
3714: waveform_sig_loopback =-8058;
3715: waveform_sig_loopback =-7936;
3716: waveform_sig_loopback =-6828;
3717: waveform_sig_loopback =-5514;
3718: waveform_sig_loopback =-7226;
3719: waveform_sig_loopback =-8418;
3720: waveform_sig_loopback =-6189;
3721: waveform_sig_loopback =-7200;
3722: waveform_sig_loopback =-6830;
3723: waveform_sig_loopback =-7488;
3724: waveform_sig_loopback =-7354;
3725: waveform_sig_loopback =-6114;
3726: waveform_sig_loopback =-7811;
3727: waveform_sig_loopback =-7140;
3728: waveform_sig_loopback =-7016;
3729: waveform_sig_loopback =-6804;
3730: waveform_sig_loopback =-8158;
3731: waveform_sig_loopback =-6137;
3732: waveform_sig_loopback =-7125;
3733: waveform_sig_loopback =-8354;
3734: waveform_sig_loopback =-6020;
3735: waveform_sig_loopback =-7317;
3736: waveform_sig_loopback =-7735;
3737: waveform_sig_loopback =-7167;
3738: waveform_sig_loopback =-6265;
3739: waveform_sig_loopback =-8058;
3740: waveform_sig_loopback =-7638;
3741: waveform_sig_loopback =-5921;
3742: waveform_sig_loopback =-7656;
3743: waveform_sig_loopback =-8240;
3744: waveform_sig_loopback =-6405;
3745: waveform_sig_loopback =-6332;
3746: waveform_sig_loopback =-8602;
3747: waveform_sig_loopback =-7510;
3748: waveform_sig_loopback =-5262;
3749: waveform_sig_loopback =-8949;
3750: waveform_sig_loopback =-5616;
3751: waveform_sig_loopback =-7723;
3752: waveform_sig_loopback =-10341;
3753: waveform_sig_loopback =-3912;
3754: waveform_sig_loopback =-7147;
3755: waveform_sig_loopback =-8173;
3756: waveform_sig_loopback =-7951;
3757: waveform_sig_loopback =-7351;
3758: waveform_sig_loopback =-5304;
3759: waveform_sig_loopback =-7733;
3760: waveform_sig_loopback =-8627;
3761: waveform_sig_loopback =-5992;
3762: waveform_sig_loopback =-7808;
3763: waveform_sig_loopback =-6652;
3764: waveform_sig_loopback =-7635;
3765: waveform_sig_loopback =-7678;
3766: waveform_sig_loopback =-5909;
3767: waveform_sig_loopback =-8159;
3768: waveform_sig_loopback =-7145;
3769: waveform_sig_loopback =-6893;
3770: waveform_sig_loopback =-7145;
3771: waveform_sig_loopback =-7940;
3772: waveform_sig_loopback =-6227;
3773: waveform_sig_loopback =-7307;
3774: waveform_sig_loopback =-8104;
3775: waveform_sig_loopback =-6165;
3776: waveform_sig_loopback =-7310;
3777: waveform_sig_loopback =-7667;
3778: waveform_sig_loopback =-7046;
3779: waveform_sig_loopback =-6302;
3780: waveform_sig_loopback =-7981;
3781: waveform_sig_loopback =-7499;
3782: waveform_sig_loopback =-5871;
3783: waveform_sig_loopback =-7522;
3784: waveform_sig_loopback =-8297;
3785: waveform_sig_loopback =-6023;
3786: waveform_sig_loopback =-6242;
3787: waveform_sig_loopback =-8746;
3788: waveform_sig_loopback =-6918;
3789: waveform_sig_loopback =-5394;
3790: waveform_sig_loopback =-8735;
3791: waveform_sig_loopback =-5047;
3792: waveform_sig_loopback =-8221;
3793: waveform_sig_loopback =-9486;
3794: waveform_sig_loopback =-3725;
3795: waveform_sig_loopback =-7253;
3796: waveform_sig_loopback =-7466;
3797: waveform_sig_loopback =-8117;
3798: waveform_sig_loopback =-6742;
3799: waveform_sig_loopback =-4920;
3800: waveform_sig_loopback =-7927;
3801: waveform_sig_loopback =-7783;
3802: waveform_sig_loopback =-5891;
3803: waveform_sig_loopback =-7529;
3804: waveform_sig_loopback =-6004;
3805: waveform_sig_loopback =-7700;
3806: waveform_sig_loopback =-6918;
3807: waveform_sig_loopback =-5581;
3808: waveform_sig_loopback =-7979;
3809: waveform_sig_loopback =-6442;
3810: waveform_sig_loopback =-6633;
3811: waveform_sig_loopback =-6717;
3812: waveform_sig_loopback =-7433;
3813: waveform_sig_loopback =-5716;
3814: waveform_sig_loopback =-6994;
3815: waveform_sig_loopback =-7441;
3816: waveform_sig_loopback =-5713;
3817: waveform_sig_loopback =-6890;
3818: waveform_sig_loopback =-6921;
3819: waveform_sig_loopback =-6701;
3820: waveform_sig_loopback =-5610;
3821: waveform_sig_loopback =-7431;
3822: waveform_sig_loopback =-7097;
3823: waveform_sig_loopback =-4935;
3824: waveform_sig_loopback =-7255;
3825: waveform_sig_loopback =-7644;
3826: waveform_sig_loopback =-5118;
3827: waveform_sig_loopback =-6107;
3828: waveform_sig_loopback =-7836;
3829: waveform_sig_loopback =-6163;
3830: waveform_sig_loopback =-5107;
3831: waveform_sig_loopback =-7665;
3832: waveform_sig_loopback =-4673;
3833: waveform_sig_loopback =-7651;
3834: waveform_sig_loopback =-8445;
3835: waveform_sig_loopback =-3421;
3836: waveform_sig_loopback =-6215;
3837: waveform_sig_loopback =-6963;
3838: waveform_sig_loopback =-7449;
3839: waveform_sig_loopback =-5656;
3840: waveform_sig_loopback =-4457;
3841: waveform_sig_loopback =-7047;
3842: waveform_sig_loopback =-7001;
3843: waveform_sig_loopback =-5190;
3844: waveform_sig_loopback =-6625;
3845: waveform_sig_loopback =-5176;
3846: waveform_sig_loopback =-7030;
3847: waveform_sig_loopback =-5899;
3848: waveform_sig_loopback =-4750;
3849: waveform_sig_loopback =-7251;
3850: waveform_sig_loopback =-5392;
3851: waveform_sig_loopback =-5848;
3852: waveform_sig_loopback =-5896;
3853: waveform_sig_loopback =-6294;
3854: waveform_sig_loopback =-5014;
3855: waveform_sig_loopback =-5993;
3856: waveform_sig_loopback =-6337;
3857: waveform_sig_loopback =-5119;
3858: waveform_sig_loopback =-5496;
3859: waveform_sig_loopback =-6299;
3860: waveform_sig_loopback =-5600;
3861: waveform_sig_loopback =-4422;
3862: waveform_sig_loopback =-6880;
3863: waveform_sig_loopback =-5578;
3864: waveform_sig_loopback =-4059;
3865: waveform_sig_loopback =-6432;
3866: waveform_sig_loopback =-6251;
3867: waveform_sig_loopback =-4252;
3868: waveform_sig_loopback =-4889;
3869: waveform_sig_loopback =-6716;
3870: waveform_sig_loopback =-5139;
3871: waveform_sig_loopback =-3913;
3872: waveform_sig_loopback =-6466;
3873: waveform_sig_loopback =-3519;
3874: waveform_sig_loopback =-6649;
3875: waveform_sig_loopback =-7027;
3876: waveform_sig_loopback =-2315;
3877: waveform_sig_loopback =-4926;
3878: waveform_sig_loopback =-6044;
3879: waveform_sig_loopback =-6043;
3880: waveform_sig_loopback =-4276;
3881: waveform_sig_loopback =-3535;
3882: waveform_sig_loopback =-5732;
3883: waveform_sig_loopback =-5672;
3884: waveform_sig_loopback =-4041;
3885: waveform_sig_loopback =-5227;
3886: waveform_sig_loopback =-4033;
3887: waveform_sig_loopback =-5800;
3888: waveform_sig_loopback =-4335;
3889: waveform_sig_loopback =-3846;
3890: waveform_sig_loopback =-5811;
3891: waveform_sig_loopback =-3858;
3892: waveform_sig_loopback =-4829;
3893: waveform_sig_loopback =-4283;
3894: waveform_sig_loopback =-5145;
3895: waveform_sig_loopback =-3652;
3896: waveform_sig_loopback =-4465;
3897: waveform_sig_loopback =-5337;
3898: waveform_sig_loopback =-3413;
3899: waveform_sig_loopback =-4227;
3900: waveform_sig_loopback =-5144;
3901: waveform_sig_loopback =-3788;
3902: waveform_sig_loopback =-3366;
3903: waveform_sig_loopback =-5424;
3904: waveform_sig_loopback =-3928;
3905: waveform_sig_loopback =-2918;
3906: waveform_sig_loopback =-4913;
3907: waveform_sig_loopback =-4714;
3908: waveform_sig_loopback =-2836;
3909: waveform_sig_loopback =-3554;
3910: waveform_sig_loopback =-5231;
3911: waveform_sig_loopback =-3649;
3912: waveform_sig_loopback =-2353;
3913: waveform_sig_loopback =-5209;
3914: waveform_sig_loopback =-1925;
3915: waveform_sig_loopback =-5229;
3916: waveform_sig_loopback =-5616;
3917: waveform_sig_loopback =-651;
3918: waveform_sig_loopback =-3502;
3919: waveform_sig_loopback =-4679;
3920: waveform_sig_loopback =-4513;
3921: waveform_sig_loopback =-2670;
3922: waveform_sig_loopback =-2043;
3923: waveform_sig_loopback =-4101;
3924: waveform_sig_loopback =-4436;
3925: waveform_sig_loopback =-2327;
3926: waveform_sig_loopback =-3484;
3927: waveform_sig_loopback =-2789;
3928: waveform_sig_loopback =-4071;
3929: waveform_sig_loopback =-2742;
3930: waveform_sig_loopback =-2333;
3931: waveform_sig_loopback =-4031;
3932: waveform_sig_loopback =-2566;
3933: waveform_sig_loopback =-3101;
3934: waveform_sig_loopback =-2654;
3935: waveform_sig_loopback =-3645;
3936: waveform_sig_loopback =-1896;
3937: waveform_sig_loopback =-3030;
3938: waveform_sig_loopback =-3572;
3939: waveform_sig_loopback =-1683;
3940: waveform_sig_loopback =-2833;
3941: waveform_sig_loopback =-3433;
3942: waveform_sig_loopback =-1908;
3943: waveform_sig_loopback =-1899;
3944: waveform_sig_loopback =-3871;
3945: waveform_sig_loopback =-2071;
3946: waveform_sig_loopback =-1329;
3947: waveform_sig_loopback =-3279;
3948: waveform_sig_loopback =-3039;
3949: waveform_sig_loopback =-1200;
3950: waveform_sig_loopback =-1667;
3951: waveform_sig_loopback =-3800;
3952: waveform_sig_loopback =-1812;
3953: waveform_sig_loopback =-470;
3954: waveform_sig_loopback =-3752;
3955: waveform_sig_loopback =14;
3956: waveform_sig_loopback =-3739;
3957: waveform_sig_loopback =-3743;
3958: waveform_sig_loopback =1427;
3959: waveform_sig_loopback =-2295;
3960: waveform_sig_loopback =-2788;
3961: waveform_sig_loopback =-2345;
3962: waveform_sig_loopback =-1291;
3963: waveform_sig_loopback =-54;
3964: waveform_sig_loopback =-2574;
3965: waveform_sig_loopback =-2431;
3966: waveform_sig_loopback =-375;
3967: waveform_sig_loopback =-2062;
3968: waveform_sig_loopback =-859;
3969: waveform_sig_loopback =-2155;
3970: waveform_sig_loopback =-1014;
3971: waveform_sig_loopback =-644;
3972: waveform_sig_loopback =-2124;
3973: waveform_sig_loopback =-749;
3974: waveform_sig_loopback =-1178;
3975: waveform_sig_loopback =-973;
3976: waveform_sig_loopback =-1897;
3977: waveform_sig_loopback =292;
3978: waveform_sig_loopback =-1484;
3979: waveform_sig_loopback =-1799;
3980: waveform_sig_loopback =487;
3981: waveform_sig_loopback =-1301;
3982: waveform_sig_loopback =-1405;
3983: waveform_sig_loopback =-25;
3984: waveform_sig_loopback =-426;
3985: waveform_sig_loopback =-1508;
3986: waveform_sig_loopback =-540;
3987: waveform_sig_loopback =513;
3988: waveform_sig_loopback =-1182;
3989: waveform_sig_loopback =-1459;
3990: waveform_sig_loopback =1118;
3991: waveform_sig_loopback =-157;
3992: waveform_sig_loopback =-2021;
3993: waveform_sig_loopback =578;
3994: waveform_sig_loopback =905;
3995: waveform_sig_loopback =-1765;
3996: waveform_sig_loopback =2076;
3997: waveform_sig_loopback =-2294;
3998: waveform_sig_loopback =-1443;
3999: waveform_sig_loopback =3160;
4000: waveform_sig_loopback =-579;
4001: waveform_sig_loopback =-636;
4002: waveform_sig_loopback =-745;
4003: waveform_sig_loopback =662;
4004: waveform_sig_loopback =2105;
4005: waveform_sig_loopback =-1012;
4006: waveform_sig_loopback =-379;
4007: waveform_sig_loopback =1489;
4008: waveform_sig_loopback =-273;
4009: waveform_sig_loopback =1286;
4010: waveform_sig_loopback =-535;
4011: waveform_sig_loopback =924;
4012: waveform_sig_loopback =1430;
4013: waveform_sig_loopback =-429;
4014: waveform_sig_loopback =1093;
4015: waveform_sig_loopback =858;
4016: waveform_sig_loopback =692;
4017: waveform_sig_loopback =220;
4018: waveform_sig_loopback =2207;
4019: waveform_sig_loopback =-12;
4020: waveform_sig_loopback =641;
4021: waveform_sig_loopback =2078;
4022: waveform_sig_loopback =515;
4023: waveform_sig_loopback =753;
4024: waveform_sig_loopback =1553;
4025: waveform_sig_loopback =1736;
4026: waveform_sig_loopback =230;
4027: waveform_sig_loopback =1287;
4028: waveform_sig_loopback =2706;
4029: waveform_sig_loopback =354;
4030: waveform_sig_loopback =510;
4031: waveform_sig_loopback =3183;
4032: waveform_sig_loopback =1401;
4033: waveform_sig_loopback =8;
4034: waveform_sig_loopback =2535;
4035: waveform_sig_loopback =2483;
4036: waveform_sig_loopback =440;
4037: waveform_sig_loopback =3853;
4038: waveform_sig_loopback =-727;
4039: waveform_sig_loopback =935;
4040: waveform_sig_loopback =4785;
4041: waveform_sig_loopback =1287;
4042: waveform_sig_loopback =1325;
4043: waveform_sig_loopback =922;
4044: waveform_sig_loopback =2801;
4045: waveform_sig_loopback =3865;
4046: waveform_sig_loopback =584;
4047: waveform_sig_loopback =1872;
4048: waveform_sig_loopback =3064;
4049: waveform_sig_loopback =1596;
4050: waveform_sig_loopback =3361;
4051: waveform_sig_loopback =961;
4052: waveform_sig_loopback =3095;
4053: waveform_sig_loopback =3158;
4054: waveform_sig_loopback =1239;
4055: waveform_sig_loopback =3245;
4056: waveform_sig_loopback =2482;
4057: waveform_sig_loopback =2472;
4058: waveform_sig_loopback =2313;
4059: waveform_sig_loopback =3705;
4060: waveform_sig_loopback =1927;
4061: waveform_sig_loopback =2573;
4062: waveform_sig_loopback =3586;
4063: waveform_sig_loopback =2607;
4064: waveform_sig_loopback =2352;
4065: waveform_sig_loopback =3370;
4066: waveform_sig_loopback =3700;
4067: waveform_sig_loopback =1728;
4068: waveform_sig_loopback =3321;
4069: waveform_sig_loopback =4471;
4070: waveform_sig_loopback =1872;
4071: waveform_sig_loopback =2585;
4072: waveform_sig_loopback =4891;
4073: waveform_sig_loopback =2972;
4074: waveform_sig_loopback =2030;
4075: waveform_sig_loopback =4240;
4076: waveform_sig_loopback =4108;
4077: waveform_sig_loopback =2419;
4078: waveform_sig_loopback =5395;
4079: waveform_sig_loopback =944;
4080: waveform_sig_loopback =2980;
4081: waveform_sig_loopback =6280;
4082: waveform_sig_loopback =3185;
4083: waveform_sig_loopback =2901;
4084: waveform_sig_loopback =2629;
4085: waveform_sig_loopback =4887;
4086: waveform_sig_loopback =5140;
4087: waveform_sig_loopback =2349;
4088: waveform_sig_loopback =3788;
4089: waveform_sig_loopback =4414;
4090: waveform_sig_loopback =3633;
4091: waveform_sig_loopback =4742;
4092: waveform_sig_loopback =2591;
4093: waveform_sig_loopback =5075;
4094: waveform_sig_loopback =4353;
4095: waveform_sig_loopback =3124;
4096: waveform_sig_loopback =4896;
4097: waveform_sig_loopback =3922;
4098: waveform_sig_loopback =4249;
4099: waveform_sig_loopback =3877;
4100: waveform_sig_loopback =5277;
4101: waveform_sig_loopback =3637;
4102: waveform_sig_loopback =4131;
4103: waveform_sig_loopback =5152;
4104: waveform_sig_loopback =4345;
4105: waveform_sig_loopback =3721;
4106: waveform_sig_loopback =5203;
4107: waveform_sig_loopback =5288;
4108: waveform_sig_loopback =3028;
4109: waveform_sig_loopback =5373;
4110: waveform_sig_loopback =5803;
4111: waveform_sig_loopback =3307;
4112: waveform_sig_loopback =4605;
4113: waveform_sig_loopback =6092;
4114: waveform_sig_loopback =4697;
4115: waveform_sig_loopback =3575;
4116: waveform_sig_loopback =5699;
4117: waveform_sig_loopback =5883;
4118: waveform_sig_loopback =3723;
4119: waveform_sig_loopback =7004;
4120: waveform_sig_loopback =2424;
4121: waveform_sig_loopback =4503;
4122: waveform_sig_loopback =7858;
4123: waveform_sig_loopback =4541;
4124: waveform_sig_loopback =4276;
4125: waveform_sig_loopback =4331;
4126: waveform_sig_loopback =6341;
4127: waveform_sig_loopback =6438;
4128: waveform_sig_loopback =3966;
4129: waveform_sig_loopback =5173;
4130: waveform_sig_loopback =5735;
4131: waveform_sig_loopback =5281;
4132: waveform_sig_loopback =5868;
4133: waveform_sig_loopback =4216;
4134: waveform_sig_loopback =6568;
4135: waveform_sig_loopback =5424;
4136: waveform_sig_loopback =4918;
4137: waveform_sig_loopback =6052;
4138: waveform_sig_loopback =5342;
4139: waveform_sig_loopback =5813;
4140: waveform_sig_loopback =4949;
4141: waveform_sig_loopback =6857;
4142: waveform_sig_loopback =4866;
4143: waveform_sig_loopback =5339;
4144: waveform_sig_loopback =6773;
4145: waveform_sig_loopback =5390;
4146: waveform_sig_loopback =5123;
4147: waveform_sig_loopback =6766;
4148: waveform_sig_loopback =6107;
4149: waveform_sig_loopback =4556;
4150: waveform_sig_loopback =6743;
4151: waveform_sig_loopback =6724;
4152: waveform_sig_loopback =4745;
4153: waveform_sig_loopback =5783;
4154: waveform_sig_loopback =7264;
4155: waveform_sig_loopback =5947;
4156: waveform_sig_loopback =4583;
4157: waveform_sig_loopback =7084;
4158: waveform_sig_loopback =6934;
4159: waveform_sig_loopback =4806;
4160: waveform_sig_loopback =8299;
4161: waveform_sig_loopback =3368;
4162: waveform_sig_loopback =5815;
4163: waveform_sig_loopback =9033;
4164: waveform_sig_loopback =5482;
4165: waveform_sig_loopback =5311;
4166: waveform_sig_loopback =5675;
4167: waveform_sig_loopback =7280;
4168: waveform_sig_loopback =7523;
4169: waveform_sig_loopback =5124;
4170: waveform_sig_loopback =6078;
4171: waveform_sig_loopback =7058;
4172: waveform_sig_loopback =6227;
4173: waveform_sig_loopback =6733;
4174: waveform_sig_loopback =5626;
4175: waveform_sig_loopback =7321;
4176: waveform_sig_loopback =6523;
4177: waveform_sig_loopback =6098;
4178: waveform_sig_loopback =6705;
4179: waveform_sig_loopback =6716;
4180: waveform_sig_loopback =6547;
4181: waveform_sig_loopback =5954;
4182: waveform_sig_loopback =8122;
4183: waveform_sig_loopback =5426;
4184: waveform_sig_loopback =6588;
4185: waveform_sig_loopback =7739;
4186: waveform_sig_loopback =6044;
4187: waveform_sig_loopback =6330;
4188: waveform_sig_loopback =7497;
4189: waveform_sig_loopback =6971;
4190: waveform_sig_loopback =5550;
4191: waveform_sig_loopback =7551;
4192: waveform_sig_loopback =7572;
4193: waveform_sig_loopback =5594;
4194: waveform_sig_loopback =6621;
4195: waveform_sig_loopback =8101;
4196: waveform_sig_loopback =6795;
4197: waveform_sig_loopback =5216;
4198: waveform_sig_loopback =8163;
4199: waveform_sig_loopback =7577;
4200: waveform_sig_loopback =5501;
4201: waveform_sig_loopback =9319;
4202: waveform_sig_loopback =3654;
4203: waveform_sig_loopback =6963;
4204: waveform_sig_loopback =9828;
4205: waveform_sig_loopback =5780;
4206: waveform_sig_loopback =6313;
4207: waveform_sig_loopback =6356;
4208: waveform_sig_loopback =7810;
4209: waveform_sig_loopback =8515;
4210: waveform_sig_loopback =5317;
4211: waveform_sig_loopback =6983;
4212: waveform_sig_loopback =7871;
4213: waveform_sig_loopback =6514;
4214: waveform_sig_loopback =7763;
4215: waveform_sig_loopback =5984;
4216: waveform_sig_loopback =7877;
4217: waveform_sig_loopback =7449;
4218: waveform_sig_loopback =6285;
4219: waveform_sig_loopback =7527;
4220: waveform_sig_loopback =7259;
4221: waveform_sig_loopback =6808;
4222: waveform_sig_loopback =6914;
4223: waveform_sig_loopback =8314;
4224: waveform_sig_loopback =5979;
4225: waveform_sig_loopback =7243;
4226: waveform_sig_loopback =8015;
4227: waveform_sig_loopback =6566;
4228: waveform_sig_loopback =6746;
4229: waveform_sig_loopback =8071;
4230: waveform_sig_loopback =7166;
4231: waveform_sig_loopback =6141;
4232: waveform_sig_loopback =7864;
4233: waveform_sig_loopback =7943;
4234: waveform_sig_loopback =6124;
4235: waveform_sig_loopback =6671;
4236: waveform_sig_loopback =8882;
4237: waveform_sig_loopback =6825;
4238: waveform_sig_loopback =5511;
4239: waveform_sig_loopback =9015;
4240: waveform_sig_loopback =7172;
4241: waveform_sig_loopback =6400;
4242: waveform_sig_loopback =9508;
4243: waveform_sig_loopback =3472;
4244: waveform_sig_loopback =8098;
4245: waveform_sig_loopback =9468;
4246: waveform_sig_loopback =6194;
4247: waveform_sig_loopback =6822;
4248: waveform_sig_loopback =6116;
4249: waveform_sig_loopback =8664;
4250: waveform_sig_loopback =8365;
4251: waveform_sig_loopback =5372;
4252: waveform_sig_loopback =7654;
4253: waveform_sig_loopback =7573;
4254: waveform_sig_loopback =6946;
4255: waveform_sig_loopback =7851;
4256: waveform_sig_loopback =5913;
4257: waveform_sig_loopback =8381;
4258: waveform_sig_loopback =7212;
4259: waveform_sig_loopback =6436;
4260: waveform_sig_loopback =7703;
4261: waveform_sig_loopback =7280;
4262: waveform_sig_loopback =6826;
4263: waveform_sig_loopback =6921;
4264: waveform_sig_loopback =8443;
4265: waveform_sig_loopback =5688;
4266: waveform_sig_loopback =7682;
4267: waveform_sig_loopback =7518;
4268: waveform_sig_loopback =6570;
4269: waveform_sig_loopback =7117;
4270: waveform_sig_loopback =7541;
4271: waveform_sig_loopback =7417;
4272: waveform_sig_loopback =5702;
4273: waveform_sig_loopback =8009;
4274: waveform_sig_loopback =8165;
4275: waveform_sig_loopback =5384;
4276: waveform_sig_loopback =7002;
4277: waveform_sig_loopback =8833;
4278: waveform_sig_loopback =6346;
4279: waveform_sig_loopback =5734;
4280: waveform_sig_loopback =8556;
4281: waveform_sig_loopback =6993;
4282: waveform_sig_loopback =6590;
4283: waveform_sig_loopback =8682;
4284: waveform_sig_loopback =3539;
4285: waveform_sig_loopback =8055;
4286: waveform_sig_loopback =8888;
4287: waveform_sig_loopback =6226;
4288: waveform_sig_loopback =6187;
4289: waveform_sig_loopback =6056;
4290: waveform_sig_loopback =8500;
4291: waveform_sig_loopback =7689;
4292: waveform_sig_loopback =5264;
4293: waveform_sig_loopback =7333;
4294: waveform_sig_loopback =7027;
4295: waveform_sig_loopback =6756;
4296: waveform_sig_loopback =7319;
4297: waveform_sig_loopback =5534;
4298: waveform_sig_loopback =8144;
4299: waveform_sig_loopback =6599;
4300: waveform_sig_loopback =6109;
4301: waveform_sig_loopback =7386;
4302: waveform_sig_loopback =6683;
4303: waveform_sig_loopback =6349;
4304: waveform_sig_loopback =6779;
4305: waveform_sig_loopback =7552;
4306: waveform_sig_loopback =5464;
4307: waveform_sig_loopback =7139;
4308: waveform_sig_loopback =6947;
4309: waveform_sig_loopback =6523;
4310: waveform_sig_loopback =5911;
4311: waveform_sig_loopback =7393;
4312: waveform_sig_loopback =6992;
4313: waveform_sig_loopback =4840;
4314: waveform_sig_loopback =7838;
4315: waveform_sig_loopback =7067;
4316: waveform_sig_loopback =4930;
4317: waveform_sig_loopback =6839;
4318: waveform_sig_loopback =7581;
4319: waveform_sig_loopback =5944;
4320: waveform_sig_loopback =5201;
4321: waveform_sig_loopback =7846;
4322: waveform_sig_loopback =6394;
4323: waveform_sig_loopback =5791;
4324: waveform_sig_loopback =8072;
4325: waveform_sig_loopback =2813;
4326: waveform_sig_loopback =7351;
4327: waveform_sig_loopback =8204;
4328: waveform_sig_loopback =5454;
4329: waveform_sig_loopback =5334;
4330: waveform_sig_loopback =5418;
4331: waveform_sig_loopback =7732;
4332: waveform_sig_loopback =6756;
4333: waveform_sig_loopback =4548;
4334: waveform_sig_loopback =6579;
4335: waveform_sig_loopback =6065;
4336: waveform_sig_loopback =6177;
4337: waveform_sig_loopback =6244;
4338: waveform_sig_loopback =4781;
4339: waveform_sig_loopback =7446;
4340: waveform_sig_loopback =5351;
4341: waveform_sig_loopback =5541;
4342: waveform_sig_loopback =6432;
4343: waveform_sig_loopback =5563;
4344: waveform_sig_loopback =5783;
4345: waveform_sig_loopback =5584;
4346: waveform_sig_loopback =6699;
4347: waveform_sig_loopback =4739;
4348: waveform_sig_loopback =5814;
4349: waveform_sig_loopback =6443;
4350: waveform_sig_loopback =5212;
4351: waveform_sig_loopback =4986;
4352: waveform_sig_loopback =6775;
4353: waveform_sig_loopback =5377;
4354: waveform_sig_loopback =4306;
4355: waveform_sig_loopback =6779;
4356: waveform_sig_loopback =5851;
4357: waveform_sig_loopback =4078;
4358: waveform_sig_loopback =5712;
4359: waveform_sig_loopback =6600;
4360: waveform_sig_loopback =4772;
4361: waveform_sig_loopback =4131;
4362: waveform_sig_loopback =6814;
4363: waveform_sig_loopback =5216;
4364: waveform_sig_loopback =4745;
4365: waveform_sig_loopback =6820;
4366: waveform_sig_loopback =1766;
4367: waveform_sig_loopback =6223;
4368: waveform_sig_loopback =7096;
4369: waveform_sig_loopback =4232;
4370: waveform_sig_loopback =3996;
4371: waveform_sig_loopback =4621;
4372: waveform_sig_loopback =6325;
4373: waveform_sig_loopback =5607;
4374: waveform_sig_loopback =3487;
4375: waveform_sig_loopback =5145;
4376: waveform_sig_loopback =5132;
4377: waveform_sig_loopback =4847;
4378: waveform_sig_loopback =4857;
4379: waveform_sig_loopback =3881;
4380: waveform_sig_loopback =5928;
4381: waveform_sig_loopback =4166;
4382: waveform_sig_loopback =4431;
4383: waveform_sig_loopback =4873;
4384: waveform_sig_loopback =4588;
4385: waveform_sig_loopback =4333;
4386: waveform_sig_loopback =4253;
4387: waveform_sig_loopback =5581;
4388: waveform_sig_loopback =3118;
4389: waveform_sig_loopback =4649;
4390: waveform_sig_loopback =5211;
4391: waveform_sig_loopback =3542;
4392: waveform_sig_loopback =3895;
4393: waveform_sig_loopback =5406;
4394: waveform_sig_loopback =3752;
4395: waveform_sig_loopback =3246;
4396: waveform_sig_loopback =5185;
4397: waveform_sig_loopback =4379;
4398: waveform_sig_loopback =2818;
4399: waveform_sig_loopback =4129;
4400: waveform_sig_loopback =5326;
4401: waveform_sig_loopback =3241;
4402: waveform_sig_loopback =2617;
4403: waveform_sig_loopback =5619;
4404: waveform_sig_loopback =3504;
4405: waveform_sig_loopback =3338;
4406: waveform_sig_loopback =5413;
4407: waveform_sig_loopback =79;
4408: waveform_sig_loopback =4988;
4409: waveform_sig_loopback =5616;
4410: waveform_sig_loopback =2443;
4411: waveform_sig_loopback =2707;
4412: waveform_sig_loopback =3141;
4413: waveform_sig_loopback =4613;
4414: waveform_sig_loopback =4346;
4415: waveform_sig_loopback =1639;
4416: waveform_sig_loopback =3738;
4417: waveform_sig_loopback =3694;
4418: waveform_sig_loopback =3015;
4419: waveform_sig_loopback =3523;
4420: waveform_sig_loopback =2239;
4421: waveform_sig_loopback =4243;
4422: waveform_sig_loopback =2756;
4423: waveform_sig_loopback =2657;
4424: waveform_sig_loopback =3288;
4425: waveform_sig_loopback =3106;
4426: waveform_sig_loopback =2447;
4427: waveform_sig_loopback =2861;
4428: waveform_sig_loopback =3918;
4429: waveform_sig_loopback =1321;
4430: waveform_sig_loopback =3254;
4431: waveform_sig_loopback =3401;
4432: waveform_sig_loopback =1775;
4433: waveform_sig_loopback =2505;
4434: waveform_sig_loopback =3519;
4435: waveform_sig_loopback =2057;
4436: waveform_sig_loopback =1750;
4437: waveform_sig_loopback =3266;
4438: waveform_sig_loopback =2893;
4439: waveform_sig_loopback =1019;
4440: waveform_sig_loopback =2385;
4441: waveform_sig_loopback =3830;
4442: waveform_sig_loopback =1175;
4443: waveform_sig_loopback =1103;
4444: waveform_sig_loopback =4062;
4445: waveform_sig_loopback =1411;
4446: waveform_sig_loopback =2036;
4447: waveform_sig_loopback =3451;
4448: waveform_sig_loopback =-1809;
4449: waveform_sig_loopback =3755;
4450: waveform_sig_loopback =3511;
4451: waveform_sig_loopback =666;
4452: waveform_sig_loopback =1173;
4453: waveform_sig_loopback =1124;
4454: waveform_sig_loopback =3158;
4455: waveform_sig_loopback =2425;
4456: waveform_sig_loopback =-362;
4457: waveform_sig_loopback =2354;
4458: waveform_sig_loopback =1553;
4459: waveform_sig_loopback =1338;
4460: waveform_sig_loopback =1813;
4461: waveform_sig_loopback =216;
4462: waveform_sig_loopback =2669;
4463: waveform_sig_loopback =865;
4464: waveform_sig_loopback =784;
4465: waveform_sig_loopback =1601;
4466: waveform_sig_loopback =1210;
4467: waveform_sig_loopback =488;
4468: waveform_sig_loopback =1399;
4469: waveform_sig_loopback =1778;
4470: waveform_sig_loopback =-532;
4471: waveform_sig_loopback =1751;
4472: waveform_sig_loopback =1137;
4473: waveform_sig_loopback =236;
4474: waveform_sig_loopback =613;
4475: waveform_sig_loopback =1500;
4476: waveform_sig_loopback =502;
4477: waveform_sig_loopback =-437;
4478: waveform_sig_loopback =1602;
4479: waveform_sig_loopback =1014;
4480: waveform_sig_loopback =-1077;
4481: waveform_sig_loopback =862;
4482: waveform_sig_loopback =1805;
4483: waveform_sig_loopback =-826;
4484: waveform_sig_loopback =-516;
4485: waveform_sig_loopback =2087;
4486: waveform_sig_loopback =-657;
4487: waveform_sig_loopback =520;
4488: waveform_sig_loopback =1212;
4489: waveform_sig_loopback =-3669;
4490: waveform_sig_loopback =2221;
4491: waveform_sig_loopback =1215;
4492: waveform_sig_loopback =-1000;
4493: waveform_sig_loopback =-799;
4494: waveform_sig_loopback =-933;
4495: waveform_sig_loopback =1754;
4496: waveform_sig_loopback =85;
4497: waveform_sig_loopback =-2159;
4498: waveform_sig_loopback =751;
4499: waveform_sig_loopback =-752;
4500: waveform_sig_loopback =-115;
4501: waveform_sig_loopback =-378;
4502: waveform_sig_loopback =-1738;
4503: waveform_sig_loopback =1110;
4504: waveform_sig_loopback =-1450;
4505: waveform_sig_loopback =-901;
4506: waveform_sig_loopback =-239;
4507: waveform_sig_loopback =-837;
4508: waveform_sig_loopback =-1262;
4509: waveform_sig_loopback =-504;
4510: waveform_sig_loopback =-295;
4511: waveform_sig_loopback =-2185;
4512: waveform_sig_loopback =-260;
4513: waveform_sig_loopback =-841;
4514: waveform_sig_loopback =-1496;
4515: waveform_sig_loopback =-1390;
4516: waveform_sig_loopback =-296;
4517: waveform_sig_loopback =-1422;
4518: waveform_sig_loopback =-2423;
4519: waveform_sig_loopback =-5;
4520: waveform_sig_loopback =-1003;
4521: waveform_sig_loopback =-3151;
4522: waveform_sig_loopback =-652;
4523: waveform_sig_loopback =-291;
4524: waveform_sig_loopback =-2777;
4525: waveform_sig_loopback =-2131;
4526: waveform_sig_loopback =-108;
4527: waveform_sig_loopback =-2377;
4528: waveform_sig_loopback =-1242;
4529: waveform_sig_loopback =-1114;
4530: waveform_sig_loopback =-5119;
4531: waveform_sig_loopback =202;
4532: waveform_sig_loopback =-738;
4533: waveform_sig_loopback =-2631;
4534: waveform_sig_loopback =-3062;
4535: waveform_sig_loopback =-2385;
4536: waveform_sig_loopback =-281;
4537: waveform_sig_loopback =-2013;
4538: waveform_sig_loopback =-3712;
4539: waveform_sig_loopback =-1342;
4540: waveform_sig_loopback =-2624;
4541: waveform_sig_loopback =-1781;
4542: waveform_sig_loopback =-2530;
4543: waveform_sig_loopback =-3326;
4544: waveform_sig_loopback =-727;
4545: waveform_sig_loopback =-3552;
4546: waveform_sig_loopback =-2450;
4547: waveform_sig_loopback =-2248;
4548: waveform_sig_loopback =-2759;
4549: waveform_sig_loopback =-2903;
4550: waveform_sig_loopback =-2465;
4551: waveform_sig_loopback =-2197;
4552: waveform_sig_loopback =-3882;
4553: waveform_sig_loopback =-2226;
4554: waveform_sig_loopback =-2494;
4555: waveform_sig_loopback =-3404;
4556: waveform_sig_loopback =-3349;
4557: waveform_sig_loopback =-1775;
4558: waveform_sig_loopback =-3556;
4559: waveform_sig_loopback =-4149;
4560: waveform_sig_loopback =-1559;
4561: waveform_sig_loopback =-3243;
4562: waveform_sig_loopback =-4611;
4563: waveform_sig_loopback =-2369;
4564: waveform_sig_loopback =-2446;
4565: waveform_sig_loopback =-4264;
4566: waveform_sig_loopback =-3998;
4567: waveform_sig_loopback =-1814;
4568: waveform_sig_loopback =-4049;
4569: waveform_sig_loopback =-3165;
4570: waveform_sig_loopback =-2820;
4571: waveform_sig_loopback =-6795;
4572: waveform_sig_loopback =-1606;
4573: waveform_sig_loopback =-2300;
4574: waveform_sig_loopback =-4672;
4575: waveform_sig_loopback =-4749;
4576: waveform_sig_loopback =-3811;
4577: waveform_sig_loopback =-2254;
4578: waveform_sig_loopback =-3627;
4579: waveform_sig_loopback =-5362;
4580: waveform_sig_loopback =-3113;
4581: waveform_sig_loopback =-4191;
4582: waveform_sig_loopback =-3494;
4583: waveform_sig_loopback =-4359;
4584: waveform_sig_loopback =-4743;
4585: waveform_sig_loopback =-2566;
4586: waveform_sig_loopback =-5268;
4587: waveform_sig_loopback =-3861;
4588: waveform_sig_loopback =-4174;
4589: waveform_sig_loopback =-4272;
4590: waveform_sig_loopback =-4515;
4591: waveform_sig_loopback =-4268;
4592: waveform_sig_loopback =-3579;
4593: waveform_sig_loopback =-5646;
4594: waveform_sig_loopback =-3902;
4595: waveform_sig_loopback =-3836;
4596: waveform_sig_loopback =-5427;
4597: waveform_sig_loopback =-4659;
4598: waveform_sig_loopback =-3356;
4599: waveform_sig_loopback =-5556;
4600: waveform_sig_loopback =-5200;
4601: waveform_sig_loopback =-3387;
4602: waveform_sig_loopback =-4861;
4603: waveform_sig_loopback =-5966;
4604: waveform_sig_loopback =-4120;
4605: waveform_sig_loopback =-3749;
4606: waveform_sig_loopback =-5916;
4607: waveform_sig_loopback =-5605;
4608: waveform_sig_loopback =-3112;
4609: waveform_sig_loopback =-5846;
4610: waveform_sig_loopback =-4481;
4611: waveform_sig_loopback =-4450;
4612: waveform_sig_loopback =-8370;
4613: waveform_sig_loopback =-2828;
4614: waveform_sig_loopback =-3946;
4615: waveform_sig_loopback =-6226;
4616: waveform_sig_loopback =-6171;
4617: waveform_sig_loopback =-5170;
4618: waveform_sig_loopback =-3992;
4619: waveform_sig_loopback =-4969;
4620: waveform_sig_loopback =-6737;
4621: waveform_sig_loopback =-4710;
4622: waveform_sig_loopback =-5530;
4623: waveform_sig_loopback =-5050;
4624: waveform_sig_loopback =-5635;
4625: waveform_sig_loopback =-5978;
4626: waveform_sig_loopback =-4498;
4627: waveform_sig_loopback =-6214;
4628: waveform_sig_loopback =-5270;
4629: waveform_sig_loopback =-5775;
4630: waveform_sig_loopback =-5256;
4631: waveform_sig_loopback =-6349;
4632: waveform_sig_loopback =-5135;
4633: waveform_sig_loopback =-5082;
4634: waveform_sig_loopback =-7311;
4635: waveform_sig_loopback =-4624;
4636: waveform_sig_loopback =-5576;
4637: waveform_sig_loopback =-6655;
4638: waveform_sig_loopback =-5856;
4639: waveform_sig_loopback =-4843;
4640: waveform_sig_loopback =-6627;
4641: waveform_sig_loopback =-6598;
4642: waveform_sig_loopback =-4645;
4643: waveform_sig_loopback =-6141;
4644: waveform_sig_loopback =-7205;
4645: waveform_sig_loopback =-5422;
4646: waveform_sig_loopback =-5014;
4647: waveform_sig_loopback =-7169;
4648: waveform_sig_loopback =-6896;
4649: waveform_sig_loopback =-4070;
4650: waveform_sig_loopback =-7429;
4651: waveform_sig_loopback =-5416;
4652: waveform_sig_loopback =-5701;
4653: waveform_sig_loopback =-9838;
4654: waveform_sig_loopback =-3441;
4655: waveform_sig_loopback =-5408;
4656: waveform_sig_loopback =-7530;
4657: waveform_sig_loopback =-6937;
4658: waveform_sig_loopback =-6613;
4659: waveform_sig_loopback =-4712;
4660: waveform_sig_loopback =-6263;
4661: waveform_sig_loopback =-8192;
4662: waveform_sig_loopback =-5243;
4663: waveform_sig_loopback =-6708;
4664: waveform_sig_loopback =-6263;
4665: waveform_sig_loopback =-6588;
4666: waveform_sig_loopback =-7152;
4667: waveform_sig_loopback =-5230;
4668: waveform_sig_loopback =-7334;
4669: waveform_sig_loopback =-6653;
4670: waveform_sig_loopback =-6298;
4671: waveform_sig_loopback =-6459;
4672: waveform_sig_loopback =-7415;
4673: waveform_sig_loopback =-5890;
4674: waveform_sig_loopback =-6353;
4675: waveform_sig_loopback =-7965;
4676: waveform_sig_loopback =-5646;
4677: waveform_sig_loopback =-6666;
4678: waveform_sig_loopback =-7363;
4679: waveform_sig_loopback =-6685;
4680: waveform_sig_loopback =-5870;
4681: waveform_sig_loopback =-7542;
4682: waveform_sig_loopback =-7320;
4683: waveform_sig_loopback =-5569;
4684: waveform_sig_loopback =-6982;
4685: waveform_sig_loopback =-8095;
4686: waveform_sig_loopback =-6127;
4687: waveform_sig_loopback =-5663;
4688: waveform_sig_loopback =-8382;
4689: waveform_sig_loopback =-7364;
4690: waveform_sig_loopback =-4774;
4691: waveform_sig_loopback =-8598;
4692: waveform_sig_loopback =-5529;
4693: waveform_sig_loopback =-7067;
4694: waveform_sig_loopback =-10328;
4695: waveform_sig_loopback =-3716;
4696: waveform_sig_loopback =-6889;
4697: waveform_sig_loopback =-7720;
4698: waveform_sig_loopback =-7808;
4699: waveform_sig_loopback =-7371;
4700: waveform_sig_loopback =-4870;
4701: waveform_sig_loopback =-7588;
4702: waveform_sig_loopback =-8428;
4703: waveform_sig_loopback =-5854;
4704: waveform_sig_loopback =-7710;
4705: waveform_sig_loopback =-6442;
4706: waveform_sig_loopback =-7567;
4707: waveform_sig_loopback =-7578;
4708: waveform_sig_loopback =-5676;
4709: waveform_sig_loopback =-8185;
4710: waveform_sig_loopback =-6951;
4711: waveform_sig_loopback =-6943;
4712: waveform_sig_loopback =-7013;
4713: waveform_sig_loopback =-7924;
4714: waveform_sig_loopback =-6324;
4715: waveform_sig_loopback =-7007;
4716: waveform_sig_loopback =-8398;
4717: waveform_sig_loopback =-5971;
4718: waveform_sig_loopback =-7442;
4719: waveform_sig_loopback =-7552;
4720: waveform_sig_loopback =-7142;
4721: waveform_sig_loopback =-6465;
4722: waveform_sig_loopback =-7658;
4723: waveform_sig_loopback =-8074;
4724: waveform_sig_loopback =-5689;
4725: waveform_sig_loopback =-7449;
4726: waveform_sig_loopback =-8805;
4727: waveform_sig_loopback =-5898;
4728: waveform_sig_loopback =-6515;
4729: waveform_sig_loopback =-8680;
4730: waveform_sig_loopback =-7268;
4731: waveform_sig_loopback =-5676;
4732: waveform_sig_loopback =-8511;
4733: waveform_sig_loopback =-5865;
4734: waveform_sig_loopback =-7793;
4735: waveform_sig_loopback =-9992;
4736: waveform_sig_loopback =-4386;
4737: waveform_sig_loopback =-6988;
4738: waveform_sig_loopback =-7792;
4739: waveform_sig_loopback =-8456;
4740: waveform_sig_loopback =-7114;
4741: waveform_sig_loopback =-5264;
4742: waveform_sig_loopback =-7856;
4743: waveform_sig_loopback =-8354;
4744: waveform_sig_loopback =-6246;
4745: waveform_sig_loopback =-7719;
4746: waveform_sig_loopback =-6473;
4747: waveform_sig_loopback =-7903;
4748: waveform_sig_loopback =-7582;
4749: waveform_sig_loopback =-5810;
4750: waveform_sig_loopback =-8341;
4751: waveform_sig_loopback =-6948;
4752: waveform_sig_loopback =-6972;
4753: waveform_sig_loopback =-7258;
4754: waveform_sig_loopback =-7707;
4755: waveform_sig_loopback =-6314;
4756: waveform_sig_loopback =-7357;
4757: waveform_sig_loopback =-7878;
4758: waveform_sig_loopback =-6385;
4759: waveform_sig_loopback =-7180;
4760: waveform_sig_loopback =-7467;
4761: waveform_sig_loopback =-7512;
4762: waveform_sig_loopback =-5800;
4763: waveform_sig_loopback =-8128;
4764: waveform_sig_loopback =-7779;
4765: waveform_sig_loopback =-5342;
4766: waveform_sig_loopback =-7895;
4767: waveform_sig_loopback =-8148;
4768: waveform_sig_loopback =-5948;
4769: waveform_sig_loopback =-6541;
4770: waveform_sig_loopback =-8259;
4771: waveform_sig_loopback =-7298;
4772: waveform_sig_loopback =-5378;
4773: waveform_sig_loopback =-8313;
4774: waveform_sig_loopback =-5731;
4775: waveform_sig_loopback =-7625;
4776: waveform_sig_loopback =-9669;
4777: waveform_sig_loopback =-4138;
4778: waveform_sig_loopback =-6706;
4779: waveform_sig_loopback =-7734;
4780: waveform_sig_loopback =-8091;
4781: waveform_sig_loopback =-6642;
4782: waveform_sig_loopback =-5194;
4783: waveform_sig_loopback =-7599;
4784: waveform_sig_loopback =-7889;
4785: waveform_sig_loopback =-6017;
4786: waveform_sig_loopback =-7353;
4787: waveform_sig_loopback =-6088;
4788: waveform_sig_loopback =-7703;
4789: waveform_sig_loopback =-6912;
4790: waveform_sig_loopback =-5600;
4791: waveform_sig_loopback =-8072;
4792: waveform_sig_loopback =-6230;
4793: waveform_sig_loopback =-6783;
4794: waveform_sig_loopback =-6812;
4795: waveform_sig_loopback =-7117;
4796: waveform_sig_loopback =-6147;
4797: waveform_sig_loopback =-6613;
4798: waveform_sig_loopback =-7544;
4799: waveform_sig_loopback =-6055;
4800: waveform_sig_loopback =-6249;
4801: waveform_sig_loopback =-7510;
4802: waveform_sig_loopback =-6572;
4803: waveform_sig_loopback =-5304;
4804: waveform_sig_loopback =-7973;
4805: waveform_sig_loopback =-6623;
4806: waveform_sig_loopback =-5190;
4807: waveform_sig_loopback =-7164;
4808: waveform_sig_loopback =-7407;
4809: waveform_sig_loopback =-5538;
4810: waveform_sig_loopback =-5710;
4811: waveform_sig_loopback =-7791;
4812: waveform_sig_loopback =-6561;
4813: waveform_sig_loopback =-4713;
4814: waveform_sig_loopback =-7741;
4815: waveform_sig_loopback =-4891;
4816: waveform_sig_loopback =-7134;
4817: waveform_sig_loopback =-8821;
4818: waveform_sig_loopback =-3434;
4819: waveform_sig_loopback =-5987;
4820: waveform_sig_loopback =-7155;
4821: waveform_sig_loopback =-7304;
4822: waveform_sig_loopback =-5674;
4823: waveform_sig_loopback =-4668;
4824: waveform_sig_loopback =-6736;
4825: waveform_sig_loopback =-7039;
4826: waveform_sig_loopback =-5409;
4827: waveform_sig_loopback =-6202;
4828: waveform_sig_loopback =-5556;
4829: waveform_sig_loopback =-6846;
4830: waveform_sig_loopback =-5717;
4831: waveform_sig_loopback =-5207;
4832: waveform_sig_loopback =-6844;
4833: waveform_sig_loopback =-5463;
4834: waveform_sig_loopback =-6090;
4835: waveform_sig_loopback =-5453;
4836: waveform_sig_loopback =-6688;
4837: waveform_sig_loopback =-4908;
4838: waveform_sig_loopback =-5696;
4839: waveform_sig_loopback =-6910;
4840: waveform_sig_loopback =-4640;
4841: waveform_sig_loopback =-5723;
4842: waveform_sig_loopback =-6452;
4843: waveform_sig_loopback =-5327;
4844: waveform_sig_loopback =-4674;
4845: waveform_sig_loopback =-6794;
4846: waveform_sig_loopback =-5536;
4847: waveform_sig_loopback =-4276;
4848: waveform_sig_loopback =-6238;
4849: waveform_sig_loopback =-6283;
4850: waveform_sig_loopback =-4478;
4851: waveform_sig_loopback =-4667;
4852: waveform_sig_loopback =-6790;
4853: waveform_sig_loopback =-5433;
4854: waveform_sig_loopback =-3422;
4855: waveform_sig_loopback =-6905;
4856: waveform_sig_loopback =-3602;
4857: waveform_sig_loopback =-6137;
4858: waveform_sig_loopback =-7703;
4859: waveform_sig_loopback =-1963;
4860: waveform_sig_loopback =-5080;
4861: waveform_sig_loopback =-6071;
4862: waveform_sig_loopback =-5764;
4863: waveform_sig_loopback =-4692;
4864: waveform_sig_loopback =-3396;
4865: waveform_sig_loopback =-5465;
4866: waveform_sig_loopback =-6071;
4867: waveform_sig_loopback =-3885;
4868: waveform_sig_loopback =-5170;
4869: waveform_sig_loopback =-4381;
4870: waveform_sig_loopback =-5341;
4871: waveform_sig_loopback =-4712;
4872: waveform_sig_loopback =-3889;
4873: waveform_sig_loopback =-5431;
4874: waveform_sig_loopback =-4406;
4875: waveform_sig_loopback =-4558;
4876: waveform_sig_loopback =-4278;
4877: waveform_sig_loopback =-5481;
4878: waveform_sig_loopback =-3271;
4879: waveform_sig_loopback =-4726;
4880: waveform_sig_loopback =-5453;
4881: waveform_sig_loopback =-3083;
4882: waveform_sig_loopback =-4613;
4883: waveform_sig_loopback =-4907;
4884: waveform_sig_loopback =-3845;
4885: waveform_sig_loopback =-3548;
4886: waveform_sig_loopback =-5187;
4887: waveform_sig_loopback =-4213;
4888: waveform_sig_loopback =-2909;
4889: waveform_sig_loopback =-4640;
4890: waveform_sig_loopback =-5049;
4891: waveform_sig_loopback =-2823;
4892: waveform_sig_loopback =-3264;
4893: waveform_sig_loopback =-5545;
4894: waveform_sig_loopback =-3609;
4895: waveform_sig_loopback =-2151;
4896: waveform_sig_loopback =-5519;
4897: waveform_sig_loopback =-1797;
4898: waveform_sig_loopback =-5051;
4899: waveform_sig_loopback =-5995;
4900: waveform_sig_loopback =-316;
4901: waveform_sig_loopback =-3872;
4902: waveform_sig_loopback =-4425;
4903: waveform_sig_loopback =-4254;
4904: waveform_sig_loopback =-3330;
4905: waveform_sig_loopback =-1514;
4906: waveform_sig_loopback =-4206;
4907: waveform_sig_loopback =-4549;
4908: waveform_sig_loopback =-2015;
4909: waveform_sig_loopback =-3944;
4910: waveform_sig_loopback =-2533;
4911: waveform_sig_loopback =-3768;
4912: waveform_sig_loopback =-3299;
4913: waveform_sig_loopback =-1987;
4914: waveform_sig_loopback =-4143;
4915: waveform_sig_loopback =-2682;
4916: waveform_sig_loopback =-2743;
4917: waveform_sig_loopback =-3025;
4918: waveform_sig_loopback =-3542;
4919: waveform_sig_loopback =-1613;
4920: waveform_sig_loopback =-3291;
4921: waveform_sig_loopback =-3479;
4922: waveform_sig_loopback =-1586;
4923: waveform_sig_loopback =-2990;
4924: waveform_sig_loopback =-3120;
4925: waveform_sig_loopback =-2252;
4926: waveform_sig_loopback =-1841;
4927: waveform_sig_loopback =-3451;
4928: waveform_sig_loopback =-2589;
4929: waveform_sig_loopback =-1121;
4930: waveform_sig_loopback =-2984;
4931: waveform_sig_loopback =-3452;
4932: waveform_sig_loopback =-863;
4933: waveform_sig_loopback =-1741;
4934: waveform_sig_loopback =-3924;
4935: waveform_sig_loopback =-1499;
4936: waveform_sig_loopback =-861;
4937: waveform_sig_loopback =-3601;
4938: waveform_sig_loopback =150;
4939: waveform_sig_loopback =-3840;
4940: waveform_sig_loopback =-3617;
4941: waveform_sig_loopback =1228;
4942: waveform_sig_loopback =-2255;
4943: waveform_sig_loopback =-2356;
4944: waveform_sig_loopback =-2788;
4945: waveform_sig_loopback =-1276;
4946: waveform_sig_loopback =339;
4947: waveform_sig_loopback =-2834;
4948: waveform_sig_loopback =-2296;
4949: waveform_sig_loopback =-374;
4950: waveform_sig_loopback =-2250;
4951: waveform_sig_loopback =-364;
4952: waveform_sig_loopback =-2530;
4953: waveform_sig_loopback =-1103;
4954: waveform_sig_loopback =-141;
4955: waveform_sig_loopback =-2619;
4956: waveform_sig_loopback =-521;
4957: waveform_sig_loopback =-1189;
4958: waveform_sig_loopback =-1172;
4959: waveform_sig_loopback =-1514;
4960: waveform_sig_loopback =-40;
4961: waveform_sig_loopback =-1429;
4962: waveform_sig_loopback =-1516;
4963: waveform_sig_loopback =42;
4964: waveform_sig_loopback =-1003;
4965: waveform_sig_loopback =-1367;
4966: waveform_sig_loopback =-365;
4967: waveform_sig_loopback =-81;
4968: waveform_sig_loopback =-1771;
4969: waveform_sig_loopback =-530;
4970: waveform_sig_loopback =785;
4971: waveform_sig_loopback =-1436;
4972: waveform_sig_loopback =-1674;
4973: waveform_sig_loopback =1469;
4974: waveform_sig_loopback =-263;
4975: waveform_sig_loopback =-1995;
4976: waveform_sig_loopback =429;
4977: waveform_sig_loopback =752;
4978: waveform_sig_loopback =-1196;
4979: waveform_sig_loopback =1569;
4980: waveform_sig_loopback =-2177;
4981: waveform_sig_loopback =-1183;
4982: waveform_sig_loopback =2698;
4983: waveform_sig_loopback =-170;
4984: waveform_sig_loopback =-673;
4985: waveform_sig_loopback =-1072;
4986: waveform_sig_loopback =1102;
4987: waveform_sig_loopback =1704;
4988: waveform_sig_loopback =-871;
4989: waveform_sig_loopback =-126;
4990: waveform_sig_loopback =1073;
4991: waveform_sig_loopback =-68;
4992: waveform_sig_loopback =1374;
4993: waveform_sig_loopback =-745;
4994: waveform_sig_loopback =1124;
4995: waveform_sig_loopback =1254;
4996: waveform_sig_loopback =-496;
4997: waveform_sig_loopback =1448;
4998: waveform_sig_loopback =507;
4999: waveform_sig_loopback =800;
5000: waveform_sig_loopback =356;
5001: waveform_sig_loopback =1875;
5002: waveform_sig_loopback =323;
5003: waveform_sig_loopback =510;
5004: waveform_sig_loopback =1842;
5005: waveform_sig_loopback =943;
5006: waveform_sig_loopback =471;
5007: waveform_sig_loopback =1406;
5008: waveform_sig_loopback =2227;
5009: waveform_sig_loopback =-214;
5010: waveform_sig_loopback =1467;
5011: waveform_sig_loopback =2795;
5012: waveform_sig_loopback =75;
5013: waveform_sig_loopback =887;
5014: waveform_sig_loopback =2808;
5015: waveform_sig_loopback =1491;
5016: waveform_sig_loopback =327;
5017: waveform_sig_loopback =2011;
5018: waveform_sig_loopback =2828;
5019: waveform_sig_loopback =471;
5020: waveform_sig_loopback =3476;
5021: waveform_sig_loopback =-115;
5022: waveform_sig_loopback =452;
5023: waveform_sig_loopback =4720;
5024: waveform_sig_loopback =1752;
5025: waveform_sig_loopback =918;
5026: waveform_sig_loopback =1129;
5027: waveform_sig_loopback =2882;
5028: waveform_sig_loopback =3481;
5029: waveform_sig_loopback =1085;
5030: waveform_sig_loopback =1602;
5031: waveform_sig_loopback =2988;
5032: waveform_sig_loopback =1866;
5033: waveform_sig_loopback =3016;
5034: waveform_sig_loopback =1154;
5035: waveform_sig_loopback =3108;
5036: waveform_sig_loopback =2944;
5037: waveform_sig_loopback =1424;
5038: waveform_sig_loopback =3259;
5039: waveform_sig_loopback =2266;
5040: waveform_sig_loopback =2781;
5041: waveform_sig_loopback =2100;
5042: waveform_sig_loopback =3591;
5043: waveform_sig_loopback =2363;
5044: waveform_sig_loopback =2088;
5045: waveform_sig_loopback =3792;
5046: waveform_sig_loopback =2810;
5047: waveform_sig_loopback =1957;
5048: waveform_sig_loopback =3728;
5049: waveform_sig_loopback =3573;
5050: waveform_sig_loopback =1583;
5051: waveform_sig_loopback =3647;
5052: waveform_sig_loopback =4078;
5053: waveform_sig_loopback =2111;
5054: waveform_sig_loopback =2682;
5055: waveform_sig_loopback =4432;
5056: waveform_sig_loopback =3530;
5057: waveform_sig_loopback =1806;
5058: waveform_sig_loopback =3927;
5059: waveform_sig_loopback =4664;
5060: waveform_sig_loopback =1916;
5061: waveform_sig_loopback =5548;
5062: waveform_sig_loopback =1327;
5063: waveform_sig_loopback =2325;
5064: waveform_sig_loopback =6625;
5065: waveform_sig_loopback =3131;
5066: waveform_sig_loopback =2719;
5067: waveform_sig_loopback =2996;
5068: waveform_sig_loopback =4524;
5069: waveform_sig_loopback =5161;
5070: waveform_sig_loopback =2767;
5071: waveform_sig_loopback =3346;
5072: waveform_sig_loopback =4695;
5073: waveform_sig_loopback =3659;
5074: waveform_sig_loopback =4498;
5075: waveform_sig_loopback =3059;
5076: waveform_sig_loopback =4765;
5077: waveform_sig_loopback =4378;
5078: waveform_sig_loopback =3439;
5079: waveform_sig_loopback =4611;
5080: waveform_sig_loopback =4018;
5081: waveform_sig_loopback =4528;
5082: waveform_sig_loopback =3457;
5083: waveform_sig_loopback =5693;
5084: waveform_sig_loopback =3675;
5085: waveform_sig_loopback =3615;
5086: waveform_sig_loopback =5794;
5087: waveform_sig_loopback =3974;
5088: waveform_sig_loopback =3761;
5089: waveform_sig_loopback =5321;
5090: waveform_sig_loopback =4806;
5091: waveform_sig_loopback =3630;
5092: waveform_sig_loopback =4990;
5093: waveform_sig_loopback =5539;
5094: waveform_sig_loopback =3806;
5095: waveform_sig_loopback =4164;
5096: waveform_sig_loopback =6163;
5097: waveform_sig_loopback =4817;
5098: waveform_sig_loopback =3317;
5099: waveform_sig_loopback =5761;
5100: waveform_sig_loopback =6000;
5101: waveform_sig_loopback =3381;
5102: waveform_sig_loopback =7184;
5103: waveform_sig_loopback =2609;
5104: waveform_sig_loopback =4005;
5105: waveform_sig_loopback =8246;
5106: waveform_sig_loopback =4441;
5107: waveform_sig_loopback =4178;
5108: waveform_sig_loopback =4665;
5109: waveform_sig_loopback =5743;
5110: waveform_sig_loopback =6882;
5111: waveform_sig_loopback =4090;
5112: waveform_sig_loopback =4608;
5113: waveform_sig_loopback =6425;
5114: waveform_sig_loopback =4781;
5115: waveform_sig_loopback =5996;
5116: waveform_sig_loopback =4565;
5117: waveform_sig_loopback =5920;
5118: waveform_sig_loopback =6032;
5119: waveform_sig_loopback =4779;
5120: waveform_sig_loopback =5824;
5121: waveform_sig_loopback =5739;
5122: waveform_sig_loopback =5547;
5123: waveform_sig_loopback =4965;
5124: waveform_sig_loopback =7066;
5125: waveform_sig_loopback =4644;
5126: waveform_sig_loopback =5483;
5127: waveform_sig_loopback =6846;
5128: waveform_sig_loopback =5137;
5129: waveform_sig_loopback =5418;
5130: waveform_sig_loopback =6572;
5131: waveform_sig_loopback =5962;
5132: waveform_sig_loopback =4909;
5133: waveform_sig_loopback =6346;
5134: waveform_sig_loopback =6819;
5135: waveform_sig_loopback =5082;
5136: waveform_sig_loopback =5192;
5137: waveform_sig_loopback =7606;
5138: waveform_sig_loopback =5987;
5139: waveform_sig_loopback =4269;
5140: waveform_sig_loopback =7447;
5141: waveform_sig_loopback =6741;
5142: waveform_sig_loopback =4777;
5143: waveform_sig_loopback =8615;
5144: waveform_sig_loopback =3068;
5145: waveform_sig_loopback =5846;
5146: waveform_sig_loopback =9213;
5147: waveform_sig_loopback =5163;
5148: waveform_sig_loopback =5818;
5149: waveform_sig_loopback =5394;
5150: waveform_sig_loopback =7080;
5151: waveform_sig_loopback =8086;
5152: waveform_sig_loopback =4589;
5153: waveform_sig_loopback =6335;
5154: waveform_sig_loopback =7266;
5155: waveform_sig_loopback =5700;
5156: waveform_sig_loopback =7406;
5157: waveform_sig_loopback =5220;
5158: waveform_sig_loopback =7216;
5159: waveform_sig_loopback =7017;
5160: waveform_sig_loopback =5560;
5161: waveform_sig_loopback =7048;
5162: waveform_sig_loopback =6726;
5163: waveform_sig_loopback =6325;
5164: waveform_sig_loopback =6209;
5165: waveform_sig_loopback =7990;
5166: waveform_sig_loopback =5377;
5167: waveform_sig_loopback =6784;
5168: waveform_sig_loopback =7473;
5169: waveform_sig_loopback =6048;
5170: waveform_sig_loopback =6607;
5171: waveform_sig_loopback =7105;
5172: waveform_sig_loopback =7197;
5173: waveform_sig_loopback =5727;
5174: waveform_sig_loopback =7034;
5175: waveform_sig_loopback =8073;
5176: waveform_sig_loopback =5454;
5177: waveform_sig_loopback =6327;
5178: waveform_sig_loopback =8659;
5179: waveform_sig_loopback =6335;
5180: waveform_sig_loopback =5438;
5181: waveform_sig_loopback =8289;
5182: waveform_sig_loopback =7143;
5183: waveform_sig_loopback =6012;
5184: waveform_sig_loopback =9079;
5185: waveform_sig_loopback =3682;
5186: waveform_sig_loopback =7179;
5187: waveform_sig_loopback =9391;
5188: waveform_sig_loopback =6160;
5189: waveform_sig_loopback =6507;
5190: waveform_sig_loopback =5779;
5191: waveform_sig_loopback =8333;
5192: waveform_sig_loopback =8332;
5193: waveform_sig_loopback =5221;
5194: waveform_sig_loopback =7309;
5195: waveform_sig_loopback =7452;
5196: waveform_sig_loopback =6671;
5197: waveform_sig_loopback =7895;
5198: waveform_sig_loopback =5633;
5199: waveform_sig_loopback =8176;
5200: waveform_sig_loopback =7326;
5201: waveform_sig_loopback =6181;
5202: waveform_sig_loopback =7749;
5203: waveform_sig_loopback =7103;
5204: waveform_sig_loopback =6788;
5205: waveform_sig_loopback =7023;
5206: waveform_sig_loopback =8206;
5207: waveform_sig_loopback =5924;
5208: waveform_sig_loopback =7555;
5209: waveform_sig_loopback =7508;
5210: waveform_sig_loopback =6982;
5211: waveform_sig_loopback =6716;
5212: waveform_sig_loopback =7529;
5213: waveform_sig_loopback =7979;
5214: waveform_sig_loopback =5502;
5215: waveform_sig_loopback =8017;
5216: waveform_sig_loopback =8293;
5217: waveform_sig_loopback =5475;
5218: waveform_sig_loopback =7273;
5219: waveform_sig_loopback =8526;
5220: waveform_sig_loopback =6785;
5221: waveform_sig_loopback =5947;
5222: waveform_sig_loopback =8313;
5223: waveform_sig_loopback =7651;
5224: waveform_sig_loopback =6317;
5225: waveform_sig_loopback =9197;
5226: waveform_sig_loopback =4006;
5227: waveform_sig_loopback =7562;
5228: waveform_sig_loopback =9511;
5229: waveform_sig_loopback =6513;
5230: waveform_sig_loopback =6539;
5231: waveform_sig_loopback =6122;
5232: waveform_sig_loopback =8723;
5233: waveform_sig_loopback =8132;
5234: waveform_sig_loopback =5611;
5235: waveform_sig_loopback =7633;
5236: waveform_sig_loopback =7256;
5237: waveform_sig_loopback =7179;
5238: waveform_sig_loopback =7779;
5239: waveform_sig_loopback =5800;
5240: waveform_sig_loopback =8591;
5241: waveform_sig_loopback =6918;
5242: waveform_sig_loopback =6525;
5243: waveform_sig_loopback =7903;
5244: waveform_sig_loopback =6833;
5245: waveform_sig_loopback =7207;
5246: waveform_sig_loopback =6873;
5247: waveform_sig_loopback =8108;
5248: waveform_sig_loopback =6293;
5249: waveform_sig_loopback =7133;
5250: waveform_sig_loopback =7783;
5251: waveform_sig_loopback =6964;
5252: waveform_sig_loopback =6393;
5253: waveform_sig_loopback =7985;
5254: waveform_sig_loopback =7510;
5255: waveform_sig_loopback =5530;
5256: waveform_sig_loopback =8213;
5257: waveform_sig_loopback =7782;
5258: waveform_sig_loopback =5596;
5259: waveform_sig_loopback =7310;
5260: waveform_sig_loopback =8201;
5261: waveform_sig_loopback =6683;
5262: waveform_sig_loopback =5809;
5263: waveform_sig_loopback =8226;
5264: waveform_sig_loopback =7545;
5265: waveform_sig_loopback =6055;
5266: waveform_sig_loopback =8927;
5267: waveform_sig_loopback =3929;
5268: waveform_sig_loopback =7351;
5269: waveform_sig_loopback =9259;
5270: waveform_sig_loopback =6311;
5271: waveform_sig_loopback =5955;
5272: waveform_sig_loopback =6300;
5273: waveform_sig_loopback =8324;
5274: waveform_sig_loopback =7632;
5275: waveform_sig_loopback =5702;
5276: waveform_sig_loopback =6952;
5277: waveform_sig_loopback =7140;
5278: waveform_sig_loopback =6978;
5279: waveform_sig_loopback =7018;
5280: waveform_sig_loopback =5879;
5281: waveform_sig_loopback =7989;
5282: waveform_sig_loopback =6451;
5283: waveform_sig_loopback =6522;
5284: waveform_sig_loopback =7086;
5285: waveform_sig_loopback =6624;
5286: waveform_sig_loopback =6835;
5287: waveform_sig_loopback =6200;
5288: waveform_sig_loopback =7945;
5289: waveform_sig_loopback =5628;
5290: waveform_sig_loopback =6627;
5291: waveform_sig_loopback =7574;
5292: waveform_sig_loopback =6130;
5293: waveform_sig_loopback =6001;
5294: waveform_sig_loopback =7677;
5295: waveform_sig_loopback =6539;
5296: waveform_sig_loopback =5281;
5297: waveform_sig_loopback =7667;
5298: waveform_sig_loopback =6965;
5299: waveform_sig_loopback =5317;
5300: waveform_sig_loopback =6558;
5301: waveform_sig_loopback =7607;
5302: waveform_sig_loopback =6238;
5303: waveform_sig_loopback =4954;
5304: waveform_sig_loopback =7783;
5305: waveform_sig_loopback =6767;
5306: waveform_sig_loopback =5326;
5307: waveform_sig_loopback =8412;
5308: waveform_sig_loopback =2997;
5309: waveform_sig_loopback =6742;
5310: waveform_sig_loopback =8750;
5311: waveform_sig_loopback =5228;
5312: waveform_sig_loopback =5293;
5313: waveform_sig_loopback =5776;
5314: waveform_sig_loopback =7163;
5315: waveform_sig_loopback =6999;
5316: waveform_sig_loopback =4837;
5317: waveform_sig_loopback =6115;
5318: waveform_sig_loopback =6613;
5319: waveform_sig_loopback =5638;
5320: waveform_sig_loopback =6367;
5321: waveform_sig_loopback =5318;
5322: waveform_sig_loopback =6785;
5323: waveform_sig_loopback =5689;
5324: waveform_sig_loopback =5590;
5325: waveform_sig_loopback =6214;
5326: waveform_sig_loopback =5932;
5327: waveform_sig_loopback =5537;
5328: waveform_sig_loopback =5470;
5329: waveform_sig_loopback =7185;
5330: waveform_sig_loopback =4302;
5331: waveform_sig_loopback =5885;
5332: waveform_sig_loopback =6666;
5333: waveform_sig_loopback =4922;
5334: waveform_sig_loopback =5280;
5335: waveform_sig_loopback =6541;
5336: waveform_sig_loopback =5372;
5337: waveform_sig_loopback =4647;
5338: waveform_sig_loopback =6358;
5339: waveform_sig_loopback =5902;
5340: waveform_sig_loopback =4427;
5341: waveform_sig_loopback =5231;
5342: waveform_sig_loopback =6805;
5343: waveform_sig_loopback =4921;
5344: waveform_sig_loopback =3740;
5345: waveform_sig_loopback =7166;
5346: waveform_sig_loopback =5098;
5347: waveform_sig_loopback =4490;
5348: waveform_sig_loopback =7347;
5349: waveform_sig_loopback =1395;
5350: waveform_sig_loopback =6197;
5351: waveform_sig_loopback =7358;
5352: waveform_sig_loopback =3891;
5353: waveform_sig_loopback =4403;
5354: waveform_sig_loopback =4349;
5355: waveform_sig_loopback =6123;
5356: waveform_sig_loopback =6107;
5357: waveform_sig_loopback =3124;
5358: waveform_sig_loopback =5174;
5359: waveform_sig_loopback =5415;
5360: waveform_sig_loopback =4370;
5361: waveform_sig_loopback =5386;
5362: waveform_sig_loopback =3677;
5363: waveform_sig_loopback =5633;
5364: waveform_sig_loopback =4732;
5365: waveform_sig_loopback =3951;
5366: waveform_sig_loopback =4919;
5367: waveform_sig_loopback =4795;
5368: waveform_sig_loopback =3997;
5369: waveform_sig_loopback =4483;
5370: waveform_sig_loopback =5548;
5371: waveform_sig_loopback =2878;
5372: waveform_sig_loopback =5025;
5373: waveform_sig_loopback =4820;
5374: waveform_sig_loopback =3655;
5375: waveform_sig_loopback =4155;
5376: waveform_sig_loopback =4917;
5377: waveform_sig_loopback =4163;
5378: waveform_sig_loopback =3117;
5379: waveform_sig_loopback =4954;
5380: waveform_sig_loopback =4746;
5381: waveform_sig_loopback =2669;
5382: waveform_sig_loopback =3949;
5383: waveform_sig_loopback =5576;
5384: waveform_sig_loopback =3148;
5385: waveform_sig_loopback =2562;
5386: waveform_sig_loopback =5801;
5387: waveform_sig_loopback =3254;
5388: waveform_sig_loopback =3524;
5389: waveform_sig_loopback =5553;
5390: waveform_sig_loopback =-259;
5391: waveform_sig_loopback =5343;
5392: waveform_sig_loopback =5360;
5393: waveform_sig_loopback =2492;
5394: waveform_sig_loopback =3085;
5395: waveform_sig_loopback =2497;
5396: waveform_sig_loopback =5111;
5397: waveform_sig_loopback =4279;
5398: waveform_sig_loopback =1369;
5399: waveform_sig_loopback =4205;
5400: waveform_sig_loopback =3294;
5401: waveform_sig_loopback =3097;
5402: waveform_sig_loopback =3814;
5403: waveform_sig_loopback =1726;
5404: waveform_sig_loopback =4586;
5405: waveform_sig_loopback =2789;
5406: waveform_sig_loopback =2379;
5407: waveform_sig_loopback =3651;
5408: waveform_sig_loopback =2891;
5409: waveform_sig_loopback =2515;
5410: waveform_sig_loopback =3040;
5411: waveform_sig_loopback =3647;
5412: waveform_sig_loopback =1518;
5413: waveform_sig_loopback =3367;
5414: waveform_sig_loopback =3062;
5415: waveform_sig_loopback =2161;
5416: waveform_sig_loopback =2404;
5417: waveform_sig_loopback =3238;
5418: waveform_sig_loopback =2600;
5419: waveform_sig_loopback =1338;
5420: waveform_sig_loopback =3341;
5421: waveform_sig_loopback =3183;
5422: waveform_sig_loopback =638;
5423: waveform_sig_loopback =2655;
5424: waveform_sig_loopback =3843;
5425: waveform_sig_loopback =1019;
5426: waveform_sig_loopback =1376;
5427: waveform_sig_loopback =3739;
5428: waveform_sig_loopback =1524;
5429: waveform_sig_loopback =2269;
5430: waveform_sig_loopback =3157;
5431: waveform_sig_loopback =-1573;
5432: waveform_sig_loopback =3621;
5433: waveform_sig_loopback =3217;
5434: waveform_sig_loopback =1278;
5435: waveform_sig_loopback =840;
5436: waveform_sig_loopback =970;
5437: waveform_sig_loopback =3577;
5438: waveform_sig_loopback =1948;
5439: waveform_sig_loopback =7;
5440: waveform_sig_loopback =2289;
5441: waveform_sig_loopback =1291;
5442: waveform_sig_loopback =1776;
5443: waveform_sig_loopback =1587;
5444: waveform_sig_loopback =102;
5445: waveform_sig_loopback =2973;
5446: waveform_sig_loopback =588;
5447: waveform_sig_loopback =909;
5448: waveform_sig_loopback =1682;
5449: waveform_sig_loopback =964;
5450: waveform_sig_loopback =860;
5451: waveform_sig_loopback =1179;
5452: waveform_sig_loopback =1669;
5453: waveform_sig_loopback =-191;
5454: waveform_sig_loopback =1452;
5455: waveform_sig_loopback =1123;
5456: waveform_sig_loopback =530;
5457: waveform_sig_loopback =260;
5458: waveform_sig_loopback =1643;
5459: waveform_sig_loopback =708;
5460: waveform_sig_loopback =-822;
5461: waveform_sig_loopback =1959;
5462: waveform_sig_loopback =927;
5463: waveform_sig_loopback =-1260;
5464: waveform_sig_loopback =1244;
5465: waveform_sig_loopback =1417;
5466: waveform_sig_loopback =-554;
5467: waveform_sig_loopback =-362;
5468: waveform_sig_loopback =1471;
5469: waveform_sig_loopback =38;
5470: waveform_sig_loopback =89;
5471: waveform_sig_loopback =1162;
5472: waveform_sig_loopback =-3082;
5473: waveform_sig_loopback =1414;
5474: waveform_sig_loopback =1691;
5475: waveform_sig_loopback =-844;
5476: waveform_sig_loopback =-1315;
5477: waveform_sig_loopback =-383;
5478: waveform_sig_loopback =1265;
5479: waveform_sig_loopback =189;
5480: waveform_sig_loopback =-1803;
5481: waveform_sig_loopback =235;
5482: waveform_sig_loopback =-464;
5483: waveform_sig_loopback =-166;
5484: waveform_sig_loopback =-443;
5485: waveform_sig_loopback =-1594;
5486: waveform_sig_loopback =1043;
5487: waveform_sig_loopback =-1483;
5488: waveform_sig_loopback =-760;
5489: waveform_sig_loopback =-243;
5490: waveform_sig_loopback =-1076;
5491: waveform_sig_loopback =-792;
5492: waveform_sig_loopback =-906;
5493: waveform_sig_loopback =-204;
5494: waveform_sig_loopback =-1796;
5495: waveform_sig_loopback =-875;
5496: waveform_sig_loopback =-250;
5497: waveform_sig_loopback =-1642;
5498: waveform_sig_loopback =-1736;
5499: waveform_sig_loopback =310;
5500: waveform_sig_loopback =-1985;
5501: waveform_sig_loopback =-2110;
5502: waveform_sig_loopback =104;
5503: waveform_sig_loopback =-1448;
5504: waveform_sig_loopback =-2604;
5505: waveform_sig_loopback =-985;
5506: waveform_sig_loopback =-363;
5507: waveform_sig_loopback =-2328;
5508: waveform_sig_loopback =-2589;
5509: waveform_sig_loopback =49;
5510: waveform_sig_loopback =-2073;
5511: waveform_sig_loopback =-1781;
5512: waveform_sig_loopback =-606;
5513: waveform_sig_loopback =-5217;
5514: waveform_sig_loopback =-214;
5515: waveform_sig_loopback =-216;
5516: waveform_sig_loopback =-2953;
5517: waveform_sig_loopback =-3008;
5518: waveform_sig_loopback =-2126;
5519: waveform_sig_loopback =-749;
5520: waveform_sig_loopback =-1710;
5521: waveform_sig_loopback =-3644;
5522: waveform_sig_loopback =-1675;
5523: waveform_sig_loopback =-2227;
5524: waveform_sig_loopback =-2077;
5525: waveform_sig_loopback =-2491;
5526: waveform_sig_loopback =-3052;
5527: waveform_sig_loopback =-1160;
5528: waveform_sig_loopback =-3351;
5529: waveform_sig_loopback =-2296;
5530: waveform_sig_loopback =-2569;
5531: waveform_sig_loopback =-2540;
5532: waveform_sig_loopback =-2867;
5533: waveform_sig_loopback =-2890;
5534: waveform_sig_loopback =-1611;
5535: waveform_sig_loopback =-4249;
5536: waveform_sig_loopback =-2318;
5537: waveform_sig_loopback =-2056;
5538: waveform_sig_loopback =-3950;
5539: waveform_sig_loopback =-2883;
5540: waveform_sig_loopback =-1958;
5541: waveform_sig_loopback =-3805;
5542: waveform_sig_loopback =-3605;
5543: waveform_sig_loopback =-2103;
5544: waveform_sig_loopback =-3001;
5545: waveform_sig_loopback =-4471;
5546: waveform_sig_loopback =-2815;
5547: waveform_sig_loopback =-2008;
5548: waveform_sig_loopback =-4315;
5549: waveform_sig_loopback =-4288;
5550: waveform_sig_loopback =-1548;
5551: waveform_sig_loopback =-4149;
5552: waveform_sig_loopback =-3342;
5553: waveform_sig_loopback =-2406;
5554: waveform_sig_loopback =-7156;
5555: waveform_sig_loopback =-1622;
5556: waveform_sig_loopback =-2062;
5557: waveform_sig_loopback =-4912;
5558: waveform_sig_loopback =-4540;
5559: waveform_sig_loopback =-3921;
5560: waveform_sig_loopback =-2507;
5561: waveform_sig_loopback =-3191;
5562: waveform_sig_loopback =-5628;
5563: waveform_sig_loopback =-3245;
5564: waveform_sig_loopback =-3763;
5565: waveform_sig_loopback =-4054;
5566: waveform_sig_loopback =-3945;
5567: waveform_sig_loopback =-4780;
5568: waveform_sig_loopback =-3014;
5569: waveform_sig_loopback =-4607;
5570: waveform_sig_loopback =-4341;
5571: waveform_sig_loopback =-4176;
5572: waveform_sig_loopback =-3839;
5573: waveform_sig_loopback =-5058;
5574: waveform_sig_loopback =-3937;
5575: waveform_sig_loopback =-3551;
5576: waveform_sig_loopback =-5997;
5577: waveform_sig_loopback =-3394;
5578: waveform_sig_loopback =-4262;
5579: waveform_sig_loopback =-5268;
5580: waveform_sig_loopback =-4470;
5581: waveform_sig_loopback =-3781;
5582: waveform_sig_loopback =-5142;
5583: waveform_sig_loopback =-5343;
5584: waveform_sig_loopback =-3616;
5585: waveform_sig_loopback =-4564;
5586: waveform_sig_loopback =-6101;
5587: waveform_sig_loopback =-4348;
5588: waveform_sig_loopback =-3489;
5589: waveform_sig_loopback =-6050;
5590: waveform_sig_loopback =-5802;
5591: waveform_sig_loopback =-2852;
5592: waveform_sig_loopback =-6135;
5593: waveform_sig_loopback =-4477;
5594: waveform_sig_loopback =-4120;
5595: waveform_sig_loopback =-8928;
5596: waveform_sig_loopback =-2502;
5597: waveform_sig_loopback =-4083;
5598: waveform_sig_loopback =-6377;
5599: waveform_sig_loopback =-5715;
5600: waveform_sig_loopback =-5776;
5601: waveform_sig_loopback =-3559;
5602: waveform_sig_loopback =-4960;
5603: waveform_sig_loopback =-7252;
5604: waveform_sig_loopback =-4174;
5605: waveform_sig_loopback =-5733;
5606: waveform_sig_loopback =-5213;
5607: waveform_sig_loopback =-5242;
5608: waveform_sig_loopback =-6458;
5609: waveform_sig_loopback =-4108;
5610: waveform_sig_loopback =-6182;
5611: waveform_sig_loopback =-5737;
5612: waveform_sig_loopback =-5166;
5613: waveform_sig_loopback =-5536;
5614: waveform_sig_loopback =-6328;
5615: waveform_sig_loopback =-5089;
5616: waveform_sig_loopback =-5163;
5617: waveform_sig_loopback =-7160;
5618: waveform_sig_loopback =-4700;
5619: waveform_sig_loopback =-5755;
5620: waveform_sig_loopback =-6355;
5621: waveform_sig_loopback =-5805;
5622: waveform_sig_loopback =-5206;
5623: waveform_sig_loopback =-6186;
5624: waveform_sig_loopback =-6820;
5625: waveform_sig_loopback =-4782;
5626: waveform_sig_loopback =-5710;
5627: waveform_sig_loopback =-7639;
5628: waveform_sig_loopback =-5179;
5629: waveform_sig_loopback =-4863;
5630: waveform_sig_loopback =-7541;
5631: waveform_sig_loopback =-6502;
5632: waveform_sig_loopback =-4319;
5633: waveform_sig_loopback =-7375;
5634: waveform_sig_loopback =-5216;
5635: waveform_sig_loopback =-5888;
5636: waveform_sig_loopback =-9658;
5637: waveform_sig_loopback =-3520;
5638: waveform_sig_loopback =-5638;
5639: waveform_sig_loopback =-6999;
5640: waveform_sig_loopback =-7193;
5641: waveform_sig_loopback =-6778;
5642: waveform_sig_loopback =-4254;
5643: waveform_sig_loopback =-6563;
5644: waveform_sig_loopback =-8002;
5645: waveform_sig_loopback =-5224;
5646: waveform_sig_loopback =-7063;
5647: waveform_sig_loopback =-5834;
5648: waveform_sig_loopback =-6697;
5649: waveform_sig_loopback =-7411;
5650: waveform_sig_loopback =-4823;
5651: waveform_sig_loopback =-7618;
5652: waveform_sig_loopback =-6507;
5653: waveform_sig_loopback =-6231;
5654: waveform_sig_loopback =-6688;
5655: waveform_sig_loopback =-7088;
5656: waveform_sig_loopback =-6025;
5657: waveform_sig_loopback =-6440;
5658: waveform_sig_loopback =-7762;
5659: waveform_sig_loopback =-5761;
5660: waveform_sig_loopback =-6786;
5661: waveform_sig_loopback =-6971;
5662: waveform_sig_loopback =-7180;
5663: waveform_sig_loopback =-5807;
5664: waveform_sig_loopback =-7060;
5665: waveform_sig_loopback =-7890;
5666: waveform_sig_loopback =-5281;
5667: waveform_sig_loopback =-7135;
5668: waveform_sig_loopback =-8162;
5669: waveform_sig_loopback =-5700;
5670: waveform_sig_loopback =-6193;
5671: waveform_sig_loopback =-8204;
5672: waveform_sig_loopback =-7096;
5673: waveform_sig_loopback =-5283;
5674: waveform_sig_loopback =-8074;
5675: waveform_sig_loopback =-5952;
5676: waveform_sig_loopback =-6958;
5677: waveform_sig_loopback =-9932;
5678: waveform_sig_loopback =-4523;
5679: waveform_sig_loopback =-6419;
5680: waveform_sig_loopback =-7529;
5681: waveform_sig_loopback =-8276;
5682: waveform_sig_loopback =-7073;
5683: waveform_sig_loopback =-5146;
5684: waveform_sig_loopback =-7408;
5685: waveform_sig_loopback =-8242;
5686: waveform_sig_loopback =-6231;
5687: waveform_sig_loopback =-7579;
5688: waveform_sig_loopback =-6245;
5689: waveform_sig_loopback =-7760;
5690: waveform_sig_loopback =-7650;
5691: waveform_sig_loopback =-5563;
5692: waveform_sig_loopback =-8350;
5693: waveform_sig_loopback =-6733;
5694: waveform_sig_loopback =-7099;
5695: waveform_sig_loopback =-7197;
5696: waveform_sig_loopback =-7440;
5697: waveform_sig_loopback =-6809;
5698: waveform_sig_loopback =-6861;
5699: waveform_sig_loopback =-8126;
5700: waveform_sig_loopback =-6504;
5701: waveform_sig_loopback =-6963;
5702: waveform_sig_loopback =-7715;
5703: waveform_sig_loopback =-7474;
5704: waveform_sig_loopback =-5928;
5705: waveform_sig_loopback =-8118;
5706: waveform_sig_loopback =-7944;
5707: waveform_sig_loopback =-5532;
5708: waveform_sig_loopback =-7770;
5709: waveform_sig_loopback =-8371;
5710: waveform_sig_loopback =-6209;
5711: waveform_sig_loopback =-6572;
5712: waveform_sig_loopback =-8260;
5713: waveform_sig_loopback =-7706;
5714: waveform_sig_loopback =-5599;
5715: waveform_sig_loopback =-8212;
5716: waveform_sig_loopback =-6351;
5717: waveform_sig_loopback =-7290;
5718: waveform_sig_loopback =-10173;
5719: waveform_sig_loopback =-4768;
5720: waveform_sig_loopback =-6448;
5721: waveform_sig_loopback =-8120;
5722: waveform_sig_loopback =-8418;
5723: waveform_sig_loopback =-6893;
5724: waveform_sig_loopback =-5701;
5725: waveform_sig_loopback =-7569;
5726: waveform_sig_loopback =-8291;
5727: waveform_sig_loopback =-6598;
5728: waveform_sig_loopback =-7374;
5729: waveform_sig_loopback =-6734;
5730: waveform_sig_loopback =-7924;
5731: waveform_sig_loopback =-7285;
5732: waveform_sig_loopback =-6191;
5733: waveform_sig_loopback =-8190;
5734: waveform_sig_loopback =-6779;
5735: waveform_sig_loopback =-7344;
5736: waveform_sig_loopback =-6950;
5737: waveform_sig_loopback =-7794;
5738: waveform_sig_loopback =-6644;
5739: waveform_sig_loopback =-6808;
5740: waveform_sig_loopback =-8356;
5741: waveform_sig_loopback =-6358;
5742: waveform_sig_loopback =-6895;
5743: waveform_sig_loopback =-7874;
5744: waveform_sig_loopback =-7232;
5745: waveform_sig_loopback =-5917;
5746: waveform_sig_loopback =-8291;
5747: waveform_sig_loopback =-7446;
5748: waveform_sig_loopback =-5627;
5749: waveform_sig_loopback =-7857;
5750: waveform_sig_loopback =-7897;
5751: waveform_sig_loopback =-6364;
5752: waveform_sig_loopback =-6313;
5753: waveform_sig_loopback =-8069;
5754: waveform_sig_loopback =-7788;
5755: waveform_sig_loopback =-4937;
5756: waveform_sig_loopback =-8449;
5757: waveform_sig_loopback =-6000;
5758: waveform_sig_loopback =-6961;
5759: waveform_sig_loopback =-10265;
5760: waveform_sig_loopback =-4035;
5761: waveform_sig_loopback =-6450;
5762: waveform_sig_loopback =-8098;
5763: waveform_sig_loopback =-7745;
5764: waveform_sig_loopback =-6832;
5765: waveform_sig_loopback =-5420;
5766: waveform_sig_loopback =-7116;
5767: waveform_sig_loopback =-8194;
5768: waveform_sig_loopback =-6086;
5769: waveform_sig_loopback =-7007;
5770: waveform_sig_loopback =-6563;
5771: waveform_sig_loopback =-7334;
5772: waveform_sig_loopback =-6971;
5773: waveform_sig_loopback =-5963;
5774: waveform_sig_loopback =-7501;
5775: waveform_sig_loopback =-6585;
5776: waveform_sig_loopback =-6899;
5777: waveform_sig_loopback =-6353;
5778: waveform_sig_loopback =-7605;
5779: waveform_sig_loopback =-5946;
5780: waveform_sig_loopback =-6420;
5781: waveform_sig_loopback =-8066;
5782: waveform_sig_loopback =-5515;
5783: waveform_sig_loopback =-6607;
5784: waveform_sig_loopback =-7480;
5785: waveform_sig_loopback =-6270;
5786: waveform_sig_loopback =-5793;
5787: waveform_sig_loopback =-7587;
5788: waveform_sig_loopback =-6704;
5789: waveform_sig_loopback =-5440;
5790: waveform_sig_loopback =-6883;
5791: waveform_sig_loopback =-7527;
5792: waveform_sig_loopback =-5744;
5793: waveform_sig_loopback =-5428;
5794: waveform_sig_loopback =-7912;
5795: waveform_sig_loopback =-6774;
5796: waveform_sig_loopback =-4311;
5797: waveform_sig_loopback =-8121;
5798: waveform_sig_loopback =-4820;
5799: waveform_sig_loopback =-6740;
5800: waveform_sig_loopback =-9418;
5801: waveform_sig_loopback =-3007;
5802: waveform_sig_loopback =-6154;
5803: waveform_sig_loopback =-7233;
5804: waveform_sig_loopback =-6885;
5805: waveform_sig_loopback =-6239;
5806: waveform_sig_loopback =-4403;
5807: waveform_sig_loopback =-6507;
5808: waveform_sig_loopback =-7552;
5809: waveform_sig_loopback =-4930;
5810: waveform_sig_loopback =-6446;
5811: waveform_sig_loopback =-5716;
5812: waveform_sig_loopback =-6323;
5813: waveform_sig_loopback =-6311;
5814: waveform_sig_loopback =-4931;
5815: waveform_sig_loopback =-6661;
5816: waveform_sig_loopback =-5923;
5817: waveform_sig_loopback =-5693;
5818: waveform_sig_loopback =-5615;
5819: waveform_sig_loopback =-6811;
5820: waveform_sig_loopback =-4613;
5821: waveform_sig_loopback =-5927;
5822: waveform_sig_loopback =-6881;
5823: waveform_sig_loopback =-4419;
5824: waveform_sig_loopback =-6062;
5825: waveform_sig_loopback =-6094;
5826: waveform_sig_loopback =-5356;
5827: waveform_sig_loopback =-4985;
5828: waveform_sig_loopback =-6315;
5829: waveform_sig_loopback =-5935;
5830: waveform_sig_loopback =-4252;
5831: waveform_sig_loopback =-5870;
5832: waveform_sig_loopback =-6761;
5833: waveform_sig_loopback =-4295;
5834: waveform_sig_loopback =-4539;
5835: waveform_sig_loopback =-7042;
5836: waveform_sig_loopback =-5261;
5837: waveform_sig_loopback =-3540;
5838: waveform_sig_loopback =-6991;
5839: waveform_sig_loopback =-3411;
5840: waveform_sig_loopback =-6200;
5841: waveform_sig_loopback =-7884;
5842: waveform_sig_loopback =-1832;
5843: waveform_sig_loopback =-5292;
5844: waveform_sig_loopback =-5826;
5845: waveform_sig_loopback =-5903;
5846: waveform_sig_loopback =-5065;
5847: waveform_sig_loopback =-2935;
5848: waveform_sig_loopback =-5710;
5849: waveform_sig_loopback =-6206;
5850: waveform_sig_loopback =-3533;
5851: waveform_sig_loopback =-5658;
5852: waveform_sig_loopback =-4051;
5853: waveform_sig_loopback =-5349;
5854: waveform_sig_loopback =-5181;
5855: waveform_sig_loopback =-3282;
5856: waveform_sig_loopback =-5834;
5857: waveform_sig_loopback =-4370;
5858: waveform_sig_loopback =-4304;
5859: waveform_sig_loopback =-4741;
5860: waveform_sig_loopback =-5028;
5861: waveform_sig_loopback =-3470;
5862: waveform_sig_loopback =-4790;
5863: waveform_sig_loopback =-5167;
5864: waveform_sig_loopback =-3411;
5865: waveform_sig_loopback =-4522;
5866: waveform_sig_loopback =-4786;
5867: waveform_sig_loopback =-4121;
5868: waveform_sig_loopback =-3429;
5869: waveform_sig_loopback =-5042;
5870: waveform_sig_loopback =-4528;
5871: waveform_sig_loopback =-2721;
5872: waveform_sig_loopback =-4528;
5873: waveform_sig_loopback =-5382;
5874: waveform_sig_loopback =-2561;
5875: waveform_sig_loopback =-3425;
5876: waveform_sig_loopback =-5602;
5877: waveform_sig_loopback =-3364;
5878: waveform_sig_loopback =-2610;
5879: waveform_sig_loopback =-5175;
5880: waveform_sig_loopback =-1839;
5881: waveform_sig_loopback =-5248;
5882: waveform_sig_loopback =-5658;
5883: waveform_sig_loopback =-704;
5884: waveform_sig_loopback =-3757;
5885: waveform_sig_loopback =-4012;
5886: waveform_sig_loopback =-4886;
5887: waveform_sig_loopback =-2941;
5888: waveform_sig_loopback =-1551;
5889: waveform_sig_loopback =-4524;
5890: waveform_sig_loopback =-4080;
5891: waveform_sig_loopback =-2421;
5892: waveform_sig_loopback =-3862;
5893: waveform_sig_loopback =-2279;
5894: waveform_sig_loopback =-4270;
5895: waveform_sig_loopback =-3004;
5896: waveform_sig_loopback =-1936;
5897: waveform_sig_loopback =-4374;
5898: waveform_sig_loopback =-2479;
5899: waveform_sig_loopback =-2988;
5900: waveform_sig_loopback =-2939;
5901: waveform_sig_loopback =-3404;
5902: waveform_sig_loopback =-1924;
5903: waveform_sig_loopback =-3144;
5904: waveform_sig_loopback =-3365;
5905: waveform_sig_loopback =-1918;
5906: waveform_sig_loopback =-2791;
5907: waveform_sig_loopback =-3018;
5908: waveform_sig_loopback =-2676;
5909: waveform_sig_loopback =-1453;
5910: waveform_sig_loopback =-3632;
5911: waveform_sig_loopback =-2811;
5912: waveform_sig_loopback =-741;
5913: waveform_sig_loopback =-3381;
5914: waveform_sig_loopback =-3267;
5915: waveform_sig_loopback =-853;
5916: waveform_sig_loopback =-2117;
5917: waveform_sig_loopback =-3380;
5918: waveform_sig_loopback =-1977;
5919: waveform_sig_loopback =-860;
5920: waveform_sig_loopback =-3157;
5921: waveform_sig_loopback =-503;
5922: waveform_sig_loopback =-3283;
5923: waveform_sig_loopback =-3862;
5924: waveform_sig_loopback =882;
5925: waveform_sig_loopback =-1664;
5926: waveform_sig_loopback =-2740;
5927: waveform_sig_loopback =-2870;
5928: waveform_sig_loopback =-997;
5929: waveform_sig_loopback =-184;
5930: waveform_sig_loopback =-2432;
5931: waveform_sig_loopback =-2357;
5932: waveform_sig_loopback =-744;
5933: waveform_sig_loopback =-1885;
5934: waveform_sig_loopback =-640;
5935: waveform_sig_loopback =-2430;
5936: waveform_sig_loopback =-1021;
5937: waveform_sig_loopback =-424;
5938: waveform_sig_loopback =-2395;
5939: waveform_sig_loopback =-582;
5940: waveform_sig_loopback =-1347;
5941: waveform_sig_loopback =-1017;
5942: waveform_sig_loopback =-1540;
5943: waveform_sig_loopback =-265;
5944: waveform_sig_loopback =-1148;
5945: waveform_sig_loopback =-1619;
5946: waveform_sig_loopback =-183;
5947: waveform_sig_loopback =-591;
5948: waveform_sig_loopback =-1645;
5949: waveform_sig_loopback =-477;
5950: waveform_sig_loopback =400;
5951: waveform_sig_loopback =-2176;
5952: waveform_sig_loopback =-274;
5953: waveform_sig_loopback =564;
5954: waveform_sig_loopback =-1479;
5955: waveform_sig_loopback =-984;
5956: waveform_sig_loopback =543;
5957: waveform_sig_loopback =95;
5958: waveform_sig_loopback =-1695;
5959: waveform_sig_loopback =-158;
5960: waveform_sig_loopback =1422;
5961: waveform_sig_loopback =-1723;
5962: waveform_sig_loopback =1652;
5963: waveform_sig_loopback =-1559;
5964: waveform_sig_loopback =-2084;
5965: waveform_sig_loopback =3183;
5966: waveform_sig_loopback =-122;
5967: waveform_sig_loopback =-941;
5968: waveform_sig_loopback =-652;
5969: waveform_sig_loopback =777;
5970: waveform_sig_loopback =1679;
5971: waveform_sig_loopback =-537;
5972: waveform_sig_loopback =-438;
5973: waveform_sig_loopback =1187;
5974: waveform_sig_loopback =60;
5975: waveform_sig_loopback =1101;
5976: waveform_sig_loopback =-399;
5977: waveform_sig_loopback =1008;
5978: waveform_sig_loopback =1187;
5979: waveform_sig_loopback =-214;
5980: waveform_sig_loopback =1250;
5981: waveform_sig_loopback =439;
5982: waveform_sig_loopback =1201;
5983: waveform_sig_loopback =-19;
5984: waveform_sig_loopback =1856;
5985: waveform_sig_loopback =872;
5986: waveform_sig_loopback =-150;
5987: waveform_sig_loopback =2281;
5988: waveform_sig_loopback =877;
5989: waveform_sig_loopback =262;
5990: waveform_sig_loopback =1958;
5991: waveform_sig_loopback =1526;
5992: waveform_sig_loopback =295;
5993: waveform_sig_loopback =1499;
5994: waveform_sig_loopback =2270;
5995: waveform_sig_loopback =787;
5996: waveform_sig_loopback =526;
5997: waveform_sig_loopback =2787;
5998: waveform_sig_loopback =1874;
5999: waveform_sig_loopback =19;
6000: waveform_sig_loopback =2115;
6001: waveform_sig_loopback =2969;
6002: waveform_sig_loopback =197;
6003: waveform_sig_loopback =3688;
6004: waveform_sig_loopback =46;
6005: waveform_sig_loopback =83;
6006: waveform_sig_loopback =5032;
6007: waveform_sig_loopback =1662;
6008: waveform_sig_loopback =789;
6009: waveform_sig_loopback =1412;
6010: waveform_sig_loopback =2542;
6011: waveform_sig_loopback =3623;
6012: waveform_sig_loopback =1220;
6013: waveform_sig_loopback =1158;
6014: waveform_sig_loopback =3518;
6015: waveform_sig_loopback =1670;
6016: waveform_sig_loopback =2737;
6017: waveform_sig_loopback =1612;
6018: waveform_sig_loopback =2788;
6019: waveform_sig_loopback =3196;
6020: waveform_sig_loopback =1502;
6021: waveform_sig_loopback =2763;
6022: waveform_sig_loopback =2778;
6023: waveform_sig_loopback =2793;
6024: waveform_sig_loopback =1637;
6025: waveform_sig_loopback =4087;
6026: waveform_sig_loopback =2158;
6027: waveform_sig_loopback =2090;
6028: waveform_sig_loopback =3988;
6029: waveform_sig_loopback =2321;
6030: waveform_sig_loopback =2598;
6031: waveform_sig_loopback =3364;
6032: waveform_sig_loopback =3392;
6033: waveform_sig_loopback =2161;
6034: waveform_sig_loopback =3191;
6035: waveform_sig_loopback =4227;
6036: waveform_sig_loopback =2341;
6037: waveform_sig_loopback =2306;
6038: waveform_sig_loopback =4725;
6039: waveform_sig_loopback =3489;
6040: waveform_sig_loopback =1638;
6041: waveform_sig_loopback =4134;
6042: waveform_sig_loopback =4583;
6043: waveform_sig_loopback =1890;
6044: waveform_sig_loopback =5656;
6045: waveform_sig_loopback =1368;
6046: waveform_sig_loopback =2170;
6047: waveform_sig_loopback =6837;
6048: waveform_sig_loopback =2988;
6049: waveform_sig_loopback =2845;
6050: waveform_sig_loopback =3077;
6051: waveform_sig_loopback =4070;
6052: waveform_sig_loopback =5647;
6053: waveform_sig_loopback =2607;
6054: waveform_sig_loopback =3154;
6055: waveform_sig_loopback =5186;
6056: waveform_sig_loopback =3007;
6057: waveform_sig_loopback =5014;
6058: waveform_sig_loopback =3028;
6059: waveform_sig_loopback =4229;
6060: waveform_sig_loopback =5112;
6061: waveform_sig_loopback =2961;
6062: waveform_sig_loopback =4673;
6063: waveform_sig_loopback =4341;
6064: waveform_sig_loopback =4048;
6065: waveform_sig_loopback =3826;
6066: waveform_sig_loopback =5517;
6067: waveform_sig_loopback =3559;
6068: waveform_sig_loopback =4036;
6069: waveform_sig_loopback =5378;
6070: waveform_sig_loopback =4075;
6071: waveform_sig_loopback =4071;
6072: waveform_sig_loopback =4926;
6073: waveform_sig_loopback =5106;
6074: waveform_sig_loopback =3614;
6075: waveform_sig_loopback =4683;
6076: waveform_sig_loopback =5898;
6077: waveform_sig_loopback =3821;
6078: waveform_sig_loopback =3850;
6079: waveform_sig_loopback =6429;
6080: waveform_sig_loopback =4787;
6081: waveform_sig_loopback =3281;
6082: waveform_sig_loopback =5958;
6083: waveform_sig_loopback =5626;
6084: waveform_sig_loopback =3690;
6085: waveform_sig_loopback =7320;
6086: waveform_sig_loopback =2325;
6087: waveform_sig_loopback =4213;
6088: waveform_sig_loopback =8030;
6089: waveform_sig_loopback =4408;
6090: waveform_sig_loopback =4625;
6091: waveform_sig_loopback =3996;
6092: waveform_sig_loopback =6089;
6093: waveform_sig_loopback =6954;
6094: waveform_sig_loopback =3638;
6095: waveform_sig_loopback =5141;
6096: waveform_sig_loopback =6081;
6097: waveform_sig_loopback =4705;
6098: waveform_sig_loopback =6459;
6099: waveform_sig_loopback =4013;
6100: waveform_sig_loopback =6161;
6101: waveform_sig_loopback =6189;
6102: waveform_sig_loopback =4309;
6103: waveform_sig_loopback =6227;
6104: waveform_sig_loopback =5500;
6105: waveform_sig_loopback =5495;
6106: waveform_sig_loopback =5214;
6107: waveform_sig_loopback =6723;
6108: waveform_sig_loopback =4873;
6109: waveform_sig_loopback =5564;
6110: waveform_sig_loopback =6434;
6111: waveform_sig_loopback =5491;
6112: waveform_sig_loopback =5427;
6113: waveform_sig_loopback =6091;
6114: waveform_sig_loopback =6616;
6115: waveform_sig_loopback =4607;
6116: waveform_sig_loopback =6154;
6117: waveform_sig_loopback =7318;
6118: waveform_sig_loopback =4605;
6119: waveform_sig_loopback =5539;
6120: waveform_sig_loopback =7538;
6121: waveform_sig_loopback =5771;
6122: waveform_sig_loopback =4764;
6123: waveform_sig_loopback =6987;
6124: waveform_sig_loopback =6847;
6125: waveform_sig_loopback =5064;
6126: waveform_sig_loopback =8222;
6127: waveform_sig_loopback =3481;
6128: waveform_sig_loopback =5724;
6129: waveform_sig_loopback =8889;
6130: waveform_sig_loopback =5708;
6131: waveform_sig_loopback =5609;
6132: waveform_sig_loopback =5101;
6133: waveform_sig_loopback =7576;
6134: waveform_sig_loopback =7618;
6135: waveform_sig_loopback =4869;
6136: waveform_sig_loopback =6436;
6137: waveform_sig_loopback =6748;
6138: waveform_sig_loopback =6197;
6139: waveform_sig_loopback =7231;
6140: waveform_sig_loopback =5047;
6141: waveform_sig_loopback =7570;
6142: waveform_sig_loopback =6721;
6143: waveform_sig_loopback =5652;
6144: waveform_sig_loopback =7252;
6145: waveform_sig_loopback =6304;
6146: waveform_sig_loopback =6686;
6147: waveform_sig_loopback =6136;
6148: waveform_sig_loopback =7675;
6149: waveform_sig_loopback =5881;
6150: waveform_sig_loopback =6460;
6151: waveform_sig_loopback =7404;
6152: waveform_sig_loopback =6513;
6153: waveform_sig_loopback =6118;
6154: waveform_sig_loopback =7208;
6155: waveform_sig_loopback =7506;
6156: waveform_sig_loopback =5250;
6157: waveform_sig_loopback =7382;
6158: waveform_sig_loopback =7995;
6159: waveform_sig_loopback =5308;
6160: waveform_sig_loopback =6748;
6161: waveform_sig_loopback =8099;
6162: waveform_sig_loopback =6638;
6163: waveform_sig_loopback =5746;
6164: waveform_sig_loopback =7587;
6165: waveform_sig_loopback =7783;
6166: waveform_sig_loopback =5769;
6167: waveform_sig_loopback =8830;
6168: waveform_sig_loopback =4372;
6169: waveform_sig_loopback =6392;
6170: waveform_sig_loopback =9643;
6171: waveform_sig_loopback =6481;
6172: waveform_sig_loopback =5947;
6173: waveform_sig_loopback =6177;
6174: waveform_sig_loopback =8164;
6175: waveform_sig_loopback =8041;
6176: waveform_sig_loopback =5805;
6177: waveform_sig_loopback =6842;
6178: waveform_sig_loopback =7545;
6179: waveform_sig_loopback =6908;
6180: waveform_sig_loopback =7525;
6181: waveform_sig_loopback =5940;
6182: waveform_sig_loopback =8057;
6183: waveform_sig_loopback =7157;
6184: waveform_sig_loopback =6447;
6185: waveform_sig_loopback =7620;
6186: waveform_sig_loopback =6922;
6187: waveform_sig_loopback =7227;
6188: waveform_sig_loopback =6590;
6189: waveform_sig_loopback =8226;
6190: waveform_sig_loopback =6362;
6191: waveform_sig_loopback =6884;
6192: waveform_sig_loopback =7983;
6193: waveform_sig_loopback =6962;
6194: waveform_sig_loopback =6386;
6195: waveform_sig_loopback =8062;
6196: waveform_sig_loopback =7593;
6197: waveform_sig_loopback =5666;
6198: waveform_sig_loopback =8097;
6199: waveform_sig_loopback =7929;
6200: waveform_sig_loopback =5959;
6201: waveform_sig_loopback =7095;
6202: waveform_sig_loopback =8236;
6203: waveform_sig_loopback =7272;
6204: waveform_sig_loopback =5776;
6205: waveform_sig_loopback =8079;
6206: waveform_sig_loopback =8149;
6207: waveform_sig_loopback =5852;
6208: waveform_sig_loopback =9431;
6209: waveform_sig_loopback =4372;
6210: waveform_sig_loopback =6756;
6211: waveform_sig_loopback =10173;
6212: waveform_sig_loopback =6363;
6213: waveform_sig_loopback =6242;
6214: waveform_sig_loopback =6658;
6215: waveform_sig_loopback =8100;
6216: waveform_sig_loopback =8467;
6217: waveform_sig_loopback =5877;
6218: waveform_sig_loopback =6979;
6219: waveform_sig_loopback =7896;
6220: waveform_sig_loopback =6931;
6221: waveform_sig_loopback =7609;
6222: waveform_sig_loopback =6226;
6223: waveform_sig_loopback =8081;
6224: waveform_sig_loopback =7254;
6225: waveform_sig_loopback =6619;
6226: waveform_sig_loopback =7522;
6227: waveform_sig_loopback =7123;
6228: waveform_sig_loopback =7278;
6229: waveform_sig_loopback =6512;
6230: waveform_sig_loopback =8465;
6231: waveform_sig_loopback =6257;
6232: waveform_sig_loopback =6817;
6233: waveform_sig_loopback =8287;
6234: waveform_sig_loopback =6536;
6235: waveform_sig_loopback =6548;
6236: waveform_sig_loopback =8198;
6237: waveform_sig_loopback =6999;
6238: waveform_sig_loopback =6098;
6239: waveform_sig_loopback =7869;
6240: waveform_sig_loopback =7692;
6241: waveform_sig_loopback =6175;
6242: waveform_sig_loopback =6586;
6243: waveform_sig_loopback =8515;
6244: waveform_sig_loopback =6985;
6245: waveform_sig_loopback =5307;
6246: waveform_sig_loopback =8508;
6247: waveform_sig_loopback =7499;
6248: waveform_sig_loopback =5758;
6249: waveform_sig_loopback =9356;
6250: waveform_sig_loopback =3690;
6251: waveform_sig_loopback =7098;
6252: waveform_sig_loopback =9709;
6253: waveform_sig_loopback =5944;
6254: waveform_sig_loopback =6275;
6255: waveform_sig_loopback =6220;
6256: waveform_sig_loopback =7899;
6257: waveform_sig_loopback =8209;
6258: waveform_sig_loopback =5411;
6259: waveform_sig_loopback =6752;
6260: waveform_sig_loopback =7605;
6261: waveform_sig_loopback =6475;
6262: waveform_sig_loopback =7292;
6263: waveform_sig_loopback =5963;
6264: waveform_sig_loopback =7505;
6265: waveform_sig_loopback =7015;
6266: waveform_sig_loopback =6206;
6267: waveform_sig_loopback =6892;
6268: waveform_sig_loopback =7098;
6269: waveform_sig_loopback =6403;
6270: waveform_sig_loopback =6273;
6271: waveform_sig_loopback =8164;
6272: waveform_sig_loopback =5149;
6273: waveform_sig_loopback =7032;
6274: waveform_sig_loopback =7407;
6275: waveform_sig_loopback =5890;
6276: waveform_sig_loopback =6478;
6277: waveform_sig_loopback =7169;
6278: waveform_sig_loopback =6799;
6279: waveform_sig_loopback =5459;
6280: waveform_sig_loopback =7173;
6281: waveform_sig_loopback =7409;
6282: waveform_sig_loopback =5214;
6283: waveform_sig_loopback =6181;
6284: waveform_sig_loopback =8024;
6285: waveform_sig_loopback =6054;
6286: waveform_sig_loopback =4844;
6287: waveform_sig_loopback =8020;
6288: waveform_sig_loopback =6522;
6289: waveform_sig_loopback =5374;
6290: waveform_sig_loopback =8629;
6291: waveform_sig_loopback =2673;
6292: waveform_sig_loopback =6910;
6293: waveform_sig_loopback =8733;
6294: waveform_sig_loopback =5050;
6295: waveform_sig_loopback =5778;
6296: waveform_sig_loopback =5229;
6297: waveform_sig_loopback =7342;
6298: waveform_sig_loopback =7488;
6299: waveform_sig_loopback =4201;
6300: waveform_sig_loopback =6479;
6301: waveform_sig_loopback =6557;
6302: waveform_sig_loopback =5553;
6303: waveform_sig_loopback =6816;
6304: waveform_sig_loopback =4710;
6305: waveform_sig_loopback =7000;
6306: waveform_sig_loopback =6123;
6307: waveform_sig_loopback =5006;
6308: waveform_sig_loopback =6487;
6309: waveform_sig_loopback =6040;
6310: waveform_sig_loopback =5296;
6311: waveform_sig_loopback =5829;
6312: waveform_sig_loopback =6831;
6313: waveform_sig_loopback =4457;
6314: waveform_sig_loopback =6218;
6315: waveform_sig_loopback =6105;
6316: waveform_sig_loopback =5323;
6317: waveform_sig_loopback =5326;
6318: waveform_sig_loopback =6208;
6319: waveform_sig_loopback =5939;
6320: waveform_sig_loopback =4244;
6321: waveform_sig_loopback =6338;
6322: waveform_sig_loopback =6396;
6323: waveform_sig_loopback =4011;
6324: waveform_sig_loopback =5351;
6325: waveform_sig_loopback =7017;
6326: waveform_sig_loopback =4697;
6327: waveform_sig_loopback =4009;
6328: waveform_sig_loopback =6993;
6329: waveform_sig_loopback =5094;
6330: waveform_sig_loopback =4772;
6331: waveform_sig_loopback =7140;
6332: waveform_sig_loopback =1538;
6333: waveform_sig_loopback =6311;
6334: waveform_sig_loopback =7013;
6335: waveform_sig_loopback =4295;
6336: waveform_sig_loopback =4504;
6337: waveform_sig_loopback =3855;
6338: waveform_sig_loopback =6764;
6339: waveform_sig_loopback =5708;
6340: waveform_sig_loopback =3162;
6341: waveform_sig_loopback =5516;
6342: waveform_sig_loopback =4840;
6343: waveform_sig_loopback =4800;
6344: waveform_sig_loopback =5367;
6345: waveform_sig_loopback =3248;
6346: waveform_sig_loopback =6239;
6347: waveform_sig_loopback =4390;
6348: waveform_sig_loopback =3967;
6349: waveform_sig_loopback =5277;
6350: waveform_sig_loopback =4369;
6351: waveform_sig_loopback =4372;
6352: waveform_sig_loopback =4346;
6353: waveform_sig_loopback =5411;
6354: waveform_sig_loopback =3313;
6355: waveform_sig_loopback =4735;
6356: waveform_sig_loopback =4817;
6357: waveform_sig_loopback =3994;
6358: waveform_sig_loopback =3848;
6359: waveform_sig_loopback =4920;
6360: waveform_sig_loopback =4600;
6361: waveform_sig_loopback =2637;
6362: waveform_sig_loopback =4952;
6363: waveform_sig_loopback =5132;
6364: waveform_sig_loopback =2325;
6365: waveform_sig_loopback =4325;
6366: waveform_sig_loopback =5098;
6367: waveform_sig_loopback =3255;
6368: waveform_sig_loopback =3168;
6369: waveform_sig_loopback =4963;
6370: waveform_sig_loopback =3804;
6371: waveform_sig_loopback =3424;
6372: waveform_sig_loopback =5324;
6373: waveform_sig_loopback =471;
6374: waveform_sig_loopback =4481;
6375: waveform_sig_loopback =5624;
6376: waveform_sig_loopback =3067;
6377: waveform_sig_loopback =2387;
6378: waveform_sig_loopback =2824;
6379: waveform_sig_loopback =5072;
6380: waveform_sig_loopback =4082;
6381: waveform_sig_loopback =1853;
6382: waveform_sig_loopback =3648;
6383: waveform_sig_loopback =3453;
6384: waveform_sig_loopback =3393;
6385: waveform_sig_loopback =3438;
6386: waveform_sig_loopback =1914;
6387: waveform_sig_loopback =4643;
6388: waveform_sig_loopback =2606;
6389: waveform_sig_loopback =2533;
6390: waveform_sig_loopback =3623;
6391: waveform_sig_loopback =2636;
6392: waveform_sig_loopback =2896;
6393: waveform_sig_loopback =2726;
6394: waveform_sig_loopback =3558;
6395: waveform_sig_loopback =1970;
6396: waveform_sig_loopback =2775;
6397: waveform_sig_loopback =3332;
6398: waveform_sig_loopback =2413;
6399: waveform_sig_loopback =1796;
6400: waveform_sig_loopback =3864;
6401: waveform_sig_loopback =2326;
6402: waveform_sig_loopback =1135;
6403: waveform_sig_loopback =3844;
6404: waveform_sig_loopback =2644;
6405: waveform_sig_loopback =1020;
6406: waveform_sig_loopback =2628;
6407: waveform_sig_loopback =3369;
6408: waveform_sig_loopback =1714;
6409: waveform_sig_loopback =991;
6410: waveform_sig_loopback =3533;
6411: waveform_sig_loopback =2147;
6412: waveform_sig_loopback =1504;
6413: waveform_sig_loopback =3574;
6414: waveform_sig_loopback =-1373;
6415: waveform_sig_loopback =2894;
6416: waveform_sig_loopback =3954;
6417: waveform_sig_loopback =930;
6418: waveform_sig_loopback =696;
6419: waveform_sig_loopback =1432;
6420: waveform_sig_loopback =2960;
6421: waveform_sig_loopback =2322;
6422: waveform_sig_loopback =157;
6423: waveform_sig_loopback =1883;
6424: waveform_sig_loopback =1733;
6425: waveform_sig_loopback =1503;
6426: waveform_sig_loopback =1545;
6427: waveform_sig_loopback =407;
6428: waveform_sig_loopback =2655;
6429: waveform_sig_loopback =627;
6430: waveform_sig_loopback =1103;
6431: waveform_sig_loopback =1483;
6432: waveform_sig_loopback =977;
6433: waveform_sig_loopback =1116;
6434: waveform_sig_loopback =583;
6435: waveform_sig_loopback =2206;
6436: waveform_sig_loopback =-208;
6437: waveform_sig_loopback =929;
6438: waveform_sig_loopback =1898;
6439: waveform_sig_loopback =-57;
6440: waveform_sig_loopback =424;
6441: waveform_sig_loopback =1923;
6442: waveform_sig_loopback =114;
6443: waveform_sig_loopback =-145;
6444: waveform_sig_loopback =1555;
6445: waveform_sig_loopback =838;
6446: waveform_sig_loopback =-695;
6447: waveform_sig_loopback =571;
6448: waveform_sig_loopback =1756;
6449: waveform_sig_loopback =-366;
6450: waveform_sig_loopback =-881;
6451: waveform_sig_loopback =1948;
6452: waveform_sig_loopback =-41;
6453: waveform_sig_loopback =-227;
6454: waveform_sig_loopback =1737;
6455: waveform_sig_loopback =-3409;
6456: waveform_sig_loopback =1245;
6457: waveform_sig_loopback =2005;
6458: waveform_sig_loopback =-1109;
6459: waveform_sig_loopback =-1093;
6460: waveform_sig_loopback =-397;
6461: waveform_sig_loopback =956;
6462: waveform_sig_loopback =567;
6463: waveform_sig_loopback =-1872;
6464: waveform_sig_loopback =-93;
6465: waveform_sig_loopback =57;
6466: waveform_sig_loopback =-607;
6467: waveform_sig_loopback =-322;
6468: waveform_sig_loopback =-1305;
6469: waveform_sig_loopback =463;
6470: waveform_sig_loopback =-944;
6471: waveform_sig_loopback =-891;
6472: waveform_sig_loopback =-663;
6473: waveform_sig_loopback =-421;
6474: waveform_sig_loopback =-1336;
6475: waveform_sig_loopback =-901;
6476: waveform_sig_loopback =329;
6477: waveform_sig_loopback =-2592;
6478: waveform_sig_loopback =-283;
6479: waveform_sig_loopback =-465;
6480: waveform_sig_loopback =-1846;
6481: waveform_sig_loopback =-1208;
6482: waveform_sig_loopback =-331;
6483: waveform_sig_loopback =-1473;
6484: waveform_sig_loopback =-2134;
6485: waveform_sig_loopback =-349;
6486: waveform_sig_loopback =-957;
6487: waveform_sig_loopback =-2683;
6488: waveform_sig_loopback =-1270;
6489: waveform_sig_loopback =-143;
6490: waveform_sig_loopback =-2306;
6491: waveform_sig_loopback =-2815;
6492: waveform_sig_loopback =272;
6493: waveform_sig_loopback =-2196;
6494: waveform_sig_loopback =-1958;
6495: waveform_sig_loopback =-89;
6496: waveform_sig_loopback =-5706;
6497: waveform_sig_loopback =-57;
6498: waveform_sig_loopback =-66;
6499: waveform_sig_loopback =-3316;
6500: waveform_sig_loopback =-2489;
6501: waveform_sig_loopback =-2629;
6502: waveform_sig_loopback =-742;
6503: waveform_sig_loopback =-1170;
6504: waveform_sig_loopback =-4193;
6505: waveform_sig_loopback =-1368;
6506: waveform_sig_loopback =-2160;
6507: waveform_sig_loopback =-2476;
6508: waveform_sig_loopback =-1790;
6509: waveform_sig_loopback =-3611;
6510: waveform_sig_loopback =-1106;
6511: waveform_sig_loopback =-2792;
6512: waveform_sig_loopback =-3029;
6513: waveform_sig_loopback =-2057;
6514: waveform_sig_loopback =-2570;
6515: waveform_sig_loopback =-3174;
6516: waveform_sig_loopback =-2456;
6517: waveform_sig_loopback =-1911;
6518: waveform_sig_loopback =-4153;
6519: waveform_sig_loopback =-2144;
6520: waveform_sig_loopback =-2473;
6521: waveform_sig_loopback =-3546;
6522: waveform_sig_loopback =-3028;
6523: waveform_sig_loopback =-2255;
6524: waveform_sig_loopback =-3276;
6525: waveform_sig_loopback =-3898;
6526: waveform_sig_loopback =-2236;
6527: waveform_sig_loopback =-2626;
6528: waveform_sig_loopback =-4710;
6529: waveform_sig_loopback =-2880;
6530: waveform_sig_loopback =-1779;
6531: waveform_sig_loopback =-4497;
6532: waveform_sig_loopback =-4143;
6533: waveform_sig_loopback =-1615;
6534: waveform_sig_loopback =-4310;
6535: waveform_sig_loopback =-3060;
6536: waveform_sig_loopback =-2421;
6537: waveform_sig_loopback =-7351;
6538: waveform_sig_loopback =-1370;
6539: waveform_sig_loopback =-2380;
6540: waveform_sig_loopback =-4619;
6541: waveform_sig_loopback =-4408;
6542: waveform_sig_loopback =-4484;
6543: waveform_sig_loopback =-1920;
6544: waveform_sig_loopback =-3494;
6545: waveform_sig_loopback =-5693;
6546: waveform_sig_loopback =-2833;
6547: waveform_sig_loopback =-4353;
6548: waveform_sig_loopback =-3690;
6549: waveform_sig_loopback =-3805;
6550: waveform_sig_loopback =-5323;
6551: waveform_sig_loopback =-2442;
6552: waveform_sig_loopback =-4926;
6553: waveform_sig_loopback =-4431;
6554: waveform_sig_loopback =-3745;
6555: waveform_sig_loopback =-4395;
6556: waveform_sig_loopback =-4629;
6557: waveform_sig_loopback =-4139;
6558: waveform_sig_loopback =-3712;
6559: waveform_sig_loopback =-5575;
6560: waveform_sig_loopback =-3803;
6561: waveform_sig_loopback =-4216;
6562: waveform_sig_loopback =-4985;
6563: waveform_sig_loopback =-4752;
6564: waveform_sig_loopback =-3781;
6565: waveform_sig_loopback =-4780;
6566: waveform_sig_loopback =-5745;
6567: waveform_sig_loopback =-3528;
6568: waveform_sig_loopback =-4313;
6569: waveform_sig_loopback =-6483;
6570: waveform_sig_loopback =-3999;
6571: waveform_sig_loopback =-3714;
6572: waveform_sig_loopback =-6087;
6573: waveform_sig_loopback =-5354;
6574: waveform_sig_loopback =-3509;
6575: waveform_sig_loopback =-5635;
6576: waveform_sig_loopback =-4515;
6577: waveform_sig_loopback =-4404;
6578: waveform_sig_loopback =-8384;
6579: waveform_sig_loopback =-3040;
6580: waveform_sig_loopback =-3911;
6581: waveform_sig_loopback =-5876;
6582: waveform_sig_loopback =-6356;
6583: waveform_sig_loopback =-5465;
6584: waveform_sig_loopback =-3445;
6585: waveform_sig_loopback =-5288;
6586: waveform_sig_loopback =-6765;
6587: waveform_sig_loopback =-4525;
6588: waveform_sig_loopback =-5751;
6589: waveform_sig_loopback =-4848;
6590: waveform_sig_loopback =-5689;
6591: waveform_sig_loopback =-6388;
6592: waveform_sig_loopback =-3920;
6593: waveform_sig_loopback =-6533;
6594: waveform_sig_loopback =-5503;
6595: waveform_sig_loopback =-5371;
6596: waveform_sig_loopback =-5663;
6597: waveform_sig_loopback =-5975;
6598: waveform_sig_loopback =-5518;
6599: waveform_sig_loopback =-5122;
6600: waveform_sig_loopback =-6832;
6601: waveform_sig_loopback =-5246;
6602: waveform_sig_loopback =-5497;
6603: waveform_sig_loopback =-6229;
6604: waveform_sig_loopback =-6331;
6605: waveform_sig_loopback =-4713;
6606: waveform_sig_loopback =-6400;
6607: waveform_sig_loopback =-7020;
6608: waveform_sig_loopback =-4461;
6609: waveform_sig_loopback =-6100;
6610: waveform_sig_loopback =-7402;
6611: waveform_sig_loopback =-5205;
6612: waveform_sig_loopback =-5250;
6613: waveform_sig_loopback =-6976;
6614: waveform_sig_loopback =-6744;
6615: waveform_sig_loopback =-4624;
6616: waveform_sig_loopback =-6779;
6617: waveform_sig_loopback =-5837;
6618: waveform_sig_loopback =-5493;
6619: waveform_sig_loopback =-9513;
6620: waveform_sig_loopback =-4266;
6621: waveform_sig_loopback =-4945;
6622: waveform_sig_loopback =-7225;
6623: waveform_sig_loopback =-7477;
6624: waveform_sig_loopback =-6353;
6625: waveform_sig_loopback =-4836;
6626: waveform_sig_loopback =-6247;
6627: waveform_sig_loopback =-7795;
6628: waveform_sig_loopback =-5860;
6629: waveform_sig_loopback =-6514;
6630: waveform_sig_loopback =-6015;
6631: waveform_sig_loopback =-6915;
6632: waveform_sig_loopback =-7111;
6633: waveform_sig_loopback =-5186;
6634: waveform_sig_loopback =-7433;
6635: waveform_sig_loopback =-6473;
6636: waveform_sig_loopback =-6587;
6637: waveform_sig_loopback =-6394;
6638: waveform_sig_loopback =-7051;
6639: waveform_sig_loopback =-6477;
6640: waveform_sig_loopback =-6014;
6641: waveform_sig_loopback =-7790;
6642: waveform_sig_loopback =-6158;
6643: waveform_sig_loopback =-6323;
6644: waveform_sig_loopback =-7325;
6645: waveform_sig_loopback =-7072;
6646: waveform_sig_loopback =-5433;
6647: waveform_sig_loopback =-7703;
6648: waveform_sig_loopback =-7439;
6649: waveform_sig_loopback =-5354;
6650: waveform_sig_loopback =-7266;
6651: waveform_sig_loopback =-7803;
6652: waveform_sig_loopback =-6301;
6653: waveform_sig_loopback =-5914;
6654: waveform_sig_loopback =-7688;
6655: waveform_sig_loopback =-7988;
6656: waveform_sig_loopback =-4888;
6657: waveform_sig_loopback =-7809;
6658: waveform_sig_loopback =-6503;
6659: waveform_sig_loopback =-6163;
6660: waveform_sig_loopback =-10640;
6661: waveform_sig_loopback =-4321;
6662: waveform_sig_loopback =-5864;
6663: waveform_sig_loopback =-8299;
6664: waveform_sig_loopback =-7692;
6665: waveform_sig_loopback =-7160;
6666: waveform_sig_loopback =-5425;
6667: waveform_sig_loopback =-7035;
6668: waveform_sig_loopback =-8452;
6669: waveform_sig_loopback =-6229;
6670: waveform_sig_loopback =-7215;
6671: waveform_sig_loopback =-6780;
6672: waveform_sig_loopback =-7399;
6673: waveform_sig_loopback =-7487;
6674: waveform_sig_loopback =-6021;
6675: waveform_sig_loopback =-7885;
6676: waveform_sig_loopback =-6966;
6677: waveform_sig_loopback =-7184;
6678: waveform_sig_loopback =-6768;
6679: waveform_sig_loopback =-7792;
6680: waveform_sig_loopback =-6853;
6681: waveform_sig_loopback =-6367;
6682: waveform_sig_loopback =-8599;
6683: waveform_sig_loopback =-6321;
6684: waveform_sig_loopback =-6811;
6685: waveform_sig_loopback =-8024;
6686: waveform_sig_loopback =-7009;
6687: waveform_sig_loopback =-6292;
6688: waveform_sig_loopback =-8029;
6689: waveform_sig_loopback =-7520;
6690: waveform_sig_loopback =-6151;
6691: waveform_sig_loopback =-7331;
6692: waveform_sig_loopback =-8285;
6693: waveform_sig_loopback =-6713;
6694: waveform_sig_loopback =-6019;
6695: waveform_sig_loopback =-8463;
6696: waveform_sig_loopback =-7933;
6697: waveform_sig_loopback =-5082;
6698: waveform_sig_loopback =-8647;
6699: waveform_sig_loopback =-6216;
6700: waveform_sig_loopback =-6827;
6701: waveform_sig_loopback =-10792;
6702: waveform_sig_loopback =-4275;
6703: waveform_sig_loopback =-6560;
6704: waveform_sig_loopback =-8248;
6705: waveform_sig_loopback =-7999;
6706: waveform_sig_loopback =-7361;
6707: waveform_sig_loopback =-5534;
6708: waveform_sig_loopback =-7225;
6709: waveform_sig_loopback =-8820;
6710: waveform_sig_loopback =-6411;
6711: waveform_sig_loopback =-7176;
6712: waveform_sig_loopback =-7023;
6713: waveform_sig_loopback =-7548;
6714: waveform_sig_loopback =-7832;
6715: waveform_sig_loopback =-5988;
6716: waveform_sig_loopback =-7703;
6717: waveform_sig_loopback =-7421;
6718: waveform_sig_loopback =-7214;
6719: waveform_sig_loopback =-6587;
6720: waveform_sig_loopback =-8122;
6721: waveform_sig_loopback =-6499;
6722: waveform_sig_loopback =-6807;
6723: waveform_sig_loopback =-8584;
6724: waveform_sig_loopback =-5795;
6725: waveform_sig_loopback =-7491;
6726: waveform_sig_loopback =-7640;
6727: waveform_sig_loopback =-6931;
6728: waveform_sig_loopback =-6494;
6729: waveform_sig_loopback =-7649;
6730: waveform_sig_loopback =-7870;
6731: waveform_sig_loopback =-5763;
6732: waveform_sig_loopback =-7244;
6733: waveform_sig_loopback =-8513;
6734: waveform_sig_loopback =-6204;
6735: waveform_sig_loopback =-6044;
6736: waveform_sig_loopback =-8441;
6737: waveform_sig_loopback =-7528;
6738: waveform_sig_loopback =-5061;
6739: waveform_sig_loopback =-8451;
6740: waveform_sig_loopback =-5844;
6741: waveform_sig_loopback =-7045;
6742: waveform_sig_loopback =-10385;
6743: waveform_sig_loopback =-3900;
6744: waveform_sig_loopback =-6585;
6745: waveform_sig_loopback =-7998;
6746: waveform_sig_loopback =-7639;
6747: waveform_sig_loopback =-7235;
6748: waveform_sig_loopback =-5061;
6749: waveform_sig_loopback =-7121;
6750: waveform_sig_loopback =-8590;
6751: waveform_sig_loopback =-5548;
6752: waveform_sig_loopback =-7467;
6753: waveform_sig_loopback =-6484;
6754: waveform_sig_loopback =-6953;
6755: waveform_sig_loopback =-7673;
6756: waveform_sig_loopback =-5332;
6757: waveform_sig_loopback =-7730;
6758: waveform_sig_loopback =-6891;
6759: waveform_sig_loopback =-6299;
6760: waveform_sig_loopback =-6880;
6761: waveform_sig_loopback =-7403;
6762: waveform_sig_loopback =-5832;
6763: waveform_sig_loopback =-6776;
6764: waveform_sig_loopback =-7625;
6765: waveform_sig_loopback =-5754;
6766: waveform_sig_loopback =-6754;
6767: waveform_sig_loopback =-7024;
6768: waveform_sig_loopback =-6761;
6769: waveform_sig_loopback =-5636;
6770: waveform_sig_loopback =-7303;
6771: waveform_sig_loopback =-7165;
6772: waveform_sig_loopback =-5183;
6773: waveform_sig_loopback =-6789;
6774: waveform_sig_loopback =-7832;
6775: waveform_sig_loopback =-5518;
6776: waveform_sig_loopback =-5451;
6777: waveform_sig_loopback =-8067;
6778: waveform_sig_loopback =-6510;
6779: waveform_sig_loopback =-4632;
6780: waveform_sig_loopback =-7939;
6781: waveform_sig_loopback =-4744;
6782: waveform_sig_loopback =-6935;
6783: waveform_sig_loopback =-9206;
6784: waveform_sig_loopback =-3196;
6785: waveform_sig_loopback =-6247;
6786: waveform_sig_loopback =-6740;
6787: waveform_sig_loopback =-7310;
6788: waveform_sig_loopback =-6270;
6789: waveform_sig_loopback =-4073;
6790: waveform_sig_loopback =-6909;
6791: waveform_sig_loopback =-7239;
6792: waveform_sig_loopback =-4975;
6793: waveform_sig_loopback =-6806;
6794: waveform_sig_loopback =-5172;
6795: waveform_sig_loopback =-6685;
6796: waveform_sig_loopback =-6452;
6797: waveform_sig_loopback =-4434;
6798: waveform_sig_loopback =-7230;
6799: waveform_sig_loopback =-5529;
6800: waveform_sig_loopback =-5758;
6801: waveform_sig_loopback =-5944;
6802: waveform_sig_loopback =-6284;
6803: waveform_sig_loopback =-5121;
6804: waveform_sig_loopback =-5754;
6805: waveform_sig_loopback =-6668;
6806: waveform_sig_loopback =-4831;
6807: waveform_sig_loopback =-5760;
6808: waveform_sig_loopback =-6085;
6809: waveform_sig_loopback =-5762;
6810: waveform_sig_loopback =-4588;
6811: waveform_sig_loopback =-6333;
6812: waveform_sig_loopback =-6252;
6813: waveform_sig_loopback =-3884;
6814: waveform_sig_loopback =-6037;
6815: waveform_sig_loopback =-6781;
6816: waveform_sig_loopback =-4093;
6817: waveform_sig_loopback =-4884;
6818: waveform_sig_loopback =-6699;
6819: waveform_sig_loopback =-5299;
6820: waveform_sig_loopback =-3894;
6821: waveform_sig_loopback =-6422;
6822: waveform_sig_loopback =-3880;
6823: waveform_sig_loopback =-6018;
6824: waveform_sig_loopback =-7571;
6825: waveform_sig_loopback =-2477;
6826: waveform_sig_loopback =-4799;
6827: waveform_sig_loopback =-5699;
6828: waveform_sig_loopback =-6415;
6829: waveform_sig_loopback =-4491;
6830: waveform_sig_loopback =-3322;
6831: waveform_sig_loopback =-5619;
6832: waveform_sig_loopback =-5803;
6833: waveform_sig_loopback =-4144;
6834: waveform_sig_loopback =-5218;
6835: waveform_sig_loopback =-4054;
6836: waveform_sig_loopback =-5608;
6837: waveform_sig_loopback =-4786;
6838: waveform_sig_loopback =-3506;
6839: waveform_sig_loopback =-5855;
6840: waveform_sig_loopback =-4137;
6841: waveform_sig_loopback =-4610;
6842: waveform_sig_loopback =-4537;
6843: waveform_sig_loopback =-4952;
6844: waveform_sig_loopback =-3821;
6845: waveform_sig_loopback =-4523;
6846: waveform_sig_loopback =-5203;
6847: waveform_sig_loopback =-3703;
6848: waveform_sig_loopback =-4143;
6849: waveform_sig_loopback =-4890;
6850: waveform_sig_loopback =-4485;
6851: waveform_sig_loopback =-2885;
6852: waveform_sig_loopback =-5466;
6853: waveform_sig_loopback =-4427;
6854: waveform_sig_loopback =-2548;
6855: waveform_sig_loopback =-5058;
6856: waveform_sig_loopback =-4807;
6857: waveform_sig_loopback =-2986;
6858: waveform_sig_loopback =-3453;
6859: waveform_sig_loopback =-5070;
6860: waveform_sig_loopback =-4226;
6861: waveform_sig_loopback =-2071;
6862: waveform_sig_loopback =-5105;
6863: waveform_sig_loopback =-2462;
6864: waveform_sig_loopback =-4387;
6865: waveform_sig_loopback =-6318;
6866: waveform_sig_loopback =-734;
6867: waveform_sig_loopback =-3255;
6868: waveform_sig_loopback =-4567;
6869: waveform_sig_loopback =-4530;
6870: waveform_sig_loopback =-3045;
6871: waveform_sig_loopback =-1947;
6872: waveform_sig_loopback =-3935;
6873: waveform_sig_loopback =-4368;
6874: waveform_sig_loopback =-2540;
6875: waveform_sig_loopback =-3543;
6876: waveform_sig_loopback =-2658;
6877: waveform_sig_loopback =-3983;
6878: waveform_sig_loopback =-3011;
6879: waveform_sig_loopback =-2224;
6880: waveform_sig_loopback =-4096;
6881: waveform_sig_loopback =-2507;
6882: waveform_sig_loopback =-3213;
6883: waveform_sig_loopback =-2672;
6884: waveform_sig_loopback =-3482;
6885: waveform_sig_loopback =-2253;
6886: waveform_sig_loopback =-2570;
6887: waveform_sig_loopback =-3932;
6888: waveform_sig_loopback =-1766;
6889: waveform_sig_loopback =-2467;
6890: waveform_sig_loopback =-3670;
6891: waveform_sig_loopback =-2051;
6892: waveform_sig_loopback =-1759;
6893: waveform_sig_loopback =-3738;
6894: waveform_sig_loopback =-2360;
6895: waveform_sig_loopback =-1350;
6896: waveform_sig_loopback =-2968;
6897: waveform_sig_loopback =-3267;
6898: waveform_sig_loopback =-1276;
6899: waveform_sig_loopback =-1562;
6900: waveform_sig_loopback =-3604;
6901: waveform_sig_loopback =-2208;
6902: waveform_sig_loopback =-382;
6903: waveform_sig_loopback =-3586;
6904: waveform_sig_loopback =-512;
6905: waveform_sig_loopback =-2810;
6906: waveform_sig_loopback =-4521;
6907: waveform_sig_loopback =1188;
6908: waveform_sig_loopback =-1631;
6909: waveform_sig_loopback =-2979;
6910: waveform_sig_loopback =-2443;
6911: waveform_sig_loopback =-1397;
6912: waveform_sig_loopback =-177;
6913: waveform_sig_loopback =-2051;
6914: waveform_sig_loopback =-2821;
6915: waveform_sig_loopback =-484;
6916: waveform_sig_loopback =-1823;
6917: waveform_sig_loopback =-1028;
6918: waveform_sig_loopback =-1958;
6919: waveform_sig_loopback =-1331;
6920: waveform_sig_loopback =-481;
6921: waveform_sig_loopback =-2030;
6922: waveform_sig_loopback =-944;
6923: waveform_sig_loopback =-1226;
6924: waveform_sig_loopback =-794;
6925: waveform_sig_loopback =-1965;
6926: waveform_sig_loopback =49;
6927: waveform_sig_loopback =-1122;
6928: waveform_sig_loopback =-2040;
6929: waveform_sig_loopback =406;
6930: waveform_sig_loopback =-1086;
6931: waveform_sig_loopback =-1552;
6932: waveform_sig_loopback =-185;
6933: waveform_sig_loopback =-164;
6934: waveform_sig_loopback =-1593;
6935: waveform_sig_loopback =-628;
6936: waveform_sig_loopback =492;
6937: waveform_sig_loopback =-997;
6938: waveform_sig_loopback =-1596;
6939: waveform_sig_loopback =775;
6940: waveform_sig_loopback =246;
6941: waveform_sig_loopback =-1966;
6942: waveform_sig_loopback =-27;
6943: waveform_sig_loopback =1378;
6944: waveform_sig_loopback =-1840;
6945: waveform_sig_loopback =1722;
6946: waveform_sig_loopback =-1334;
6947: waveform_sig_loopback =-2444;
6948: waveform_sig_loopback =3316;
6949: waveform_sig_loopback =-151;
6950: waveform_sig_loopback =-950;
6951: waveform_sig_loopback =-466;
6952: waveform_sig_loopback =178;
6953: waveform_sig_loopback =2158;
6954: waveform_sig_loopback =-477;
6955: waveform_sig_loopback =-1002;
6956: waveform_sig_loopback =1805;
6957: waveform_sig_loopback =-411;
6958: waveform_sig_loopback =1235;
6959: waveform_sig_loopback =-168;
6960: waveform_sig_loopback =360;
6961: waveform_sig_loopback =1752;
6962: waveform_sig_loopback =-413;
6963: waveform_sig_loopback =955;
6964: waveform_sig_loopback =896;
6965: waveform_sig_loopback =789;
6966: waveform_sig_loopback =131;
6967: waveform_sig_loopback =2010;
6968: waveform_sig_loopback =439;
6969: waveform_sig_loopback =188;
6970: waveform_sig_loopback =2189;
6971: waveform_sig_loopback =643;
6972: waveform_sig_loopback =575;
6973: waveform_sig_loopback =1593;
6974: waveform_sig_loopback =1700;
6975: waveform_sig_loopback =381;
6976: waveform_sig_loopback =1140;
6977: waveform_sig_loopback =2510;
6978: waveform_sig_loopback =906;
6979: waveform_sig_loopback =83;
6980: waveform_sig_loopback =2988;
6981: waveform_sig_loopback =1965;
6982: waveform_sig_loopback =-228;
6983: waveform_sig_loopback =2333;
6984: waveform_sig_loopback =2806;
6985: waveform_sig_loopback =206;
6986: waveform_sig_loopback =3870;
6987: waveform_sig_loopback =-131;
6988: waveform_sig_loopback =101;
6989: waveform_sig_loopback =5021;
6990: waveform_sig_loopback =1436;
6991: waveform_sig_loopback =1353;
6992: waveform_sig_loopback =949;
6993: waveform_sig_loopback =2417;
6994: waveform_sig_loopback =4072;
6995: waveform_sig_loopback =848;
6996: waveform_sig_loopback =1451;
6997: waveform_sig_loopback =3333;
6998: waveform_sig_loopback =1424;
6999: waveform_sig_loopback =3339;
7000: waveform_sig_loopback =1235;
7001: waveform_sig_loopback =2609;
7002: waveform_sig_loopback =3544;
7003: waveform_sig_loopback =1135;
7004: waveform_sig_loopback =3087;
7005: waveform_sig_loopback =2626;
7006: waveform_sig_loopback =2589;
7007: waveform_sig_loopback =2083;
7008: waveform_sig_loopback =3804;
7009: waveform_sig_loopback =2079;
7010: waveform_sig_loopback =2380;
7011: waveform_sig_loopback =3734;
7012: waveform_sig_loopback =2537;
7013: waveform_sig_loopback =2546;
7014: waveform_sig_loopback =3095;
7015: waveform_sig_loopback =3902;
7016: waveform_sig_loopback =1955;
7017: waveform_sig_loopback =2867;
7018: waveform_sig_loopback =4673;
7019: waveform_sig_loopback =2208;
7020: waveform_sig_loopback =2268;
7021: waveform_sig_loopback =4814;
7022: waveform_sig_loopback =3305;
7023: waveform_sig_loopback =1957;
7024: waveform_sig_loopback =4007;
7025: waveform_sig_loopback =4447;
7026: waveform_sig_loopback =2302;
7027: waveform_sig_loopback =5280;
7028: waveform_sig_loopback =1460;
7029: waveform_sig_loopback =2315;
7030: waveform_sig_loopback =6588;
7031: waveform_sig_loopback =3238;
7032: waveform_sig_loopback =2807;
7033: waveform_sig_loopback =2591;
7034: waveform_sig_loopback =4736;
7035: waveform_sig_loopback =5371;
7036: waveform_sig_loopback =2465;
7037: waveform_sig_loopback =3560;
7038: waveform_sig_loopback =4640;
7039: waveform_sig_loopback =3467;
7040: waveform_sig_loopback =5008;
7041: waveform_sig_loopback =2659;
7042: waveform_sig_loopback =4722;
7043: waveform_sig_loopback =4737;
7044: waveform_sig_loopback =3049;
7045: waveform_sig_loopback =4967;
7046: waveform_sig_loopback =3875;
7047: waveform_sig_loopback =4363;
7048: waveform_sig_loopback =3794;
7049: waveform_sig_loopback =5387;
7050: waveform_sig_loopback =3844;
7051: waveform_sig_loopback =3821;
7052: waveform_sig_loopback =5305;
7053: waveform_sig_loopback =4460;
7054: waveform_sig_loopback =3741;
7055: waveform_sig_loopback =4821;
7056: waveform_sig_loopback =5628;
7057: waveform_sig_loopback =3224;
7058: waveform_sig_loopback =4650;
7059: waveform_sig_loopback =6028;
7060: waveform_sig_loopback =3763;
7061: waveform_sig_loopback =4233;
7062: waveform_sig_loopback =5853;
7063: waveform_sig_loopback =4791;
7064: waveform_sig_loopback =3949;
7065: waveform_sig_loopback =5327;
7066: waveform_sig_loopback =5955;
7067: waveform_sig_loopback =3668;
7068: waveform_sig_loopback =6995;
7069: waveform_sig_loopback =3073;
7070: waveform_sig_loopback =3471;
7071: waveform_sig_loopback =8051;
7072: waveform_sig_loopback =4989;
7073: waveform_sig_loopback =4091;
7074: waveform_sig_loopback =4159;
7075: waveform_sig_loopback =6177;
7076: waveform_sig_loopback =6713;
7077: waveform_sig_loopback =4193;
7078: waveform_sig_loopback =4673;
7079: waveform_sig_loopback =6021;
7080: waveform_sig_loopback =5259;
7081: waveform_sig_loopback =5957;
7082: waveform_sig_loopback =4252;
7083: waveform_sig_loopback =6231;
7084: waveform_sig_loopback =5963;
7085: waveform_sig_loopback =4639;
7086: waveform_sig_loopback =5996;
7087: waveform_sig_loopback =5428;
7088: waveform_sig_loopback =5866;
7089: waveform_sig_loopback =4871;
7090: waveform_sig_loopback =6732;
7091: waveform_sig_loopback =5240;
7092: waveform_sig_loopback =5116;
7093: waveform_sig_loopback =6643;
7094: waveform_sig_loopback =5626;
7095: waveform_sig_loopback =5049;
7096: waveform_sig_loopback =6419;
7097: waveform_sig_loopback =6466;
7098: waveform_sig_loopback =4457;
7099: waveform_sig_loopback =6434;
7100: waveform_sig_loopback =6903;
7101: waveform_sig_loopback =4860;
7102: waveform_sig_loopback =5560;
7103: waveform_sig_loopback =7098;
7104: waveform_sig_loopback =6254;
7105: waveform_sig_loopback =4587;
7106: waveform_sig_loopback =6641;
7107: waveform_sig_loopback =7410;
7108: waveform_sig_loopback =4521;
7109: waveform_sig_loopback =8287;
7110: waveform_sig_loopback =3983;
7111: waveform_sig_loopback =4840;
7112: waveform_sig_loopback =9437;
7113: waveform_sig_loopback =5656;
7114: waveform_sig_loopback =5265;
7115: waveform_sig_loopback =5707;
7116: waveform_sig_loopback =6946;
7117: waveform_sig_loopback =7860;
7118: waveform_sig_loopback =5248;
7119: waveform_sig_loopback =5805;
7120: waveform_sig_loopback =7343;
7121: waveform_sig_loopback =5917;
7122: waveform_sig_loopback =7102;
7123: waveform_sig_loopback =5519;
7124: waveform_sig_loopback =7046;
7125: waveform_sig_loopback =7029;
7126: waveform_sig_loopback =5667;
7127: waveform_sig_loopback =7025;
7128: waveform_sig_loopback =6523;
7129: waveform_sig_loopback =6715;
7130: waveform_sig_loopback =5834;
7131: waveform_sig_loopback =7842;
7132: waveform_sig_loopback =6075;
7133: waveform_sig_loopback =5983;
7134: waveform_sig_loopback =7837;
7135: waveform_sig_loopback =6275;
7136: waveform_sig_loopback =6096;
7137: waveform_sig_loopback =7551;
7138: waveform_sig_loopback =6936;
7139: waveform_sig_loopback =5759;
7140: waveform_sig_loopback =7188;
7141: waveform_sig_loopback =7640;
7142: waveform_sig_loopback =6057;
7143: waveform_sig_loopback =6049;
7144: waveform_sig_loopback =8174;
7145: waveform_sig_loopback =6991;
7146: waveform_sig_loopback =5131;
7147: waveform_sig_loopback =8033;
7148: waveform_sig_loopback =7655;
7149: waveform_sig_loopback =5539;
7150: waveform_sig_loopback =9241;
7151: waveform_sig_loopback =4192;
7152: waveform_sig_loopback =6168;
7153: waveform_sig_loopback =9964;
7154: waveform_sig_loopback =6210;
7155: waveform_sig_loopback =6222;
7156: waveform_sig_loopback =6178;
7157: waveform_sig_loopback =7818;
7158: waveform_sig_loopback =8548;
7159: waveform_sig_loopback =5639;
7160: waveform_sig_loopback =6680;
7161: waveform_sig_loopback =7936;
7162: waveform_sig_loopback =6565;
7163: waveform_sig_loopback =7758;
7164: waveform_sig_loopback =6025;
7165: waveform_sig_loopback =7712;
7166: waveform_sig_loopback =7564;
7167: waveform_sig_loopback =6256;
7168: waveform_sig_loopback =7413;
7169: waveform_sig_loopback =7276;
7170: waveform_sig_loopback =7062;
7171: waveform_sig_loopback =6400;
7172: waveform_sig_loopback =8650;
7173: waveform_sig_loopback =6006;
7174: waveform_sig_loopback =7004;
7175: waveform_sig_loopback =8164;
7176: waveform_sig_loopback =6553;
7177: waveform_sig_loopback =6961;
7178: waveform_sig_loopback =7532;
7179: waveform_sig_loopback =7723;
7180: waveform_sig_loopback =6094;
7181: waveform_sig_loopback =7415;
7182: waveform_sig_loopback =8415;
7183: waveform_sig_loopback =6030;
7184: waveform_sig_loopback =6654;
7185: waveform_sig_loopback =8735;
7186: waveform_sig_loopback =7037;
7187: waveform_sig_loopback =5712;
7188: waveform_sig_loopback =8354;
7189: waveform_sig_loopback =7823;
7190: waveform_sig_loopback =6028;
7191: waveform_sig_loopback =9444;
7192: waveform_sig_loopback =4185;
7193: waveform_sig_loopback =6901;
7194: waveform_sig_loopback =10007;
7195: waveform_sig_loopback =6364;
7196: waveform_sig_loopback =6570;
7197: waveform_sig_loopback =6211;
7198: waveform_sig_loopback =8205;
7199: waveform_sig_loopback =8659;
7200: waveform_sig_loopback =5597;
7201: waveform_sig_loopback =7080;
7202: waveform_sig_loopback =7914;
7203: waveform_sig_loopback =6650;
7204: waveform_sig_loopback =8025;
7205: waveform_sig_loopback =5946;
7206: waveform_sig_loopback =7910;
7207: waveform_sig_loopback =7769;
7208: waveform_sig_loopback =6116;
7209: waveform_sig_loopback =7701;
7210: waveform_sig_loopback =7359;
7211: waveform_sig_loopback =6793;
7212: waveform_sig_loopback =6954;
7213: waveform_sig_loopback =8270;
7214: waveform_sig_loopback =6055;
7215: waveform_sig_loopback =7292;
7216: waveform_sig_loopback =7638;
7217: waveform_sig_loopback =7014;
7218: waveform_sig_loopback =6599;
7219: waveform_sig_loopback =7547;
7220: waveform_sig_loopback =7876;
7221: waveform_sig_loopback =5590;
7222: waveform_sig_loopback =7752;
7223: waveform_sig_loopback =8105;
7224: waveform_sig_loopback =5828;
7225: waveform_sig_loopback =6788;
7226: waveform_sig_loopback =8397;
7227: waveform_sig_loopback =6924;
7228: waveform_sig_loopback =5520;
7229: waveform_sig_loopback =8313;
7230: waveform_sig_loopback =7464;
7231: waveform_sig_loopback =5962;
7232: waveform_sig_loopback =9296;
7233: waveform_sig_loopback =3691;
7234: waveform_sig_loopback =7144;
7235: waveform_sig_loopback =9496;
7236: waveform_sig_loopback =6144;
7237: waveform_sig_loopback =6419;
7238: waveform_sig_loopback =5708;
7239: waveform_sig_loopback =8332;
7240: waveform_sig_loopback =8096;
7241: waveform_sig_loopback =5216;
7242: waveform_sig_loopback =7180;
7243: waveform_sig_loopback =7121;
7244: waveform_sig_loopback =6656;
7245: waveform_sig_loopback =7573;
7246: waveform_sig_loopback =5346;
7247: waveform_sig_loopback =8050;
7248: waveform_sig_loopback =6886;
7249: waveform_sig_loopback =5887;
7250: waveform_sig_loopback =7455;
7251: waveform_sig_loopback =6540;
7252: waveform_sig_loopback =6707;
7253: waveform_sig_loopback =6335;
7254: waveform_sig_loopback =7731;
7255: waveform_sig_loopback =5854;
7256: waveform_sig_loopback =6554;
7257: waveform_sig_loopback =7335;
7258: waveform_sig_loopback =6409;
7259: waveform_sig_loopback =5975;
7260: waveform_sig_loopback =7202;
7261: waveform_sig_loopback =7138;
7262: waveform_sig_loopback =5103;
7263: waveform_sig_loopback =7261;
7264: waveform_sig_loopback =7459;
7265: waveform_sig_loopback =5100;
7266: waveform_sig_loopback =6391;
7267: waveform_sig_loopback =7778;
7268: waveform_sig_loopback =6057;
7269: waveform_sig_loopback =5238;
7270: waveform_sig_loopback =7525;
7271: waveform_sig_loopback =6735;
7272: waveform_sig_loopback =5555;
7273: waveform_sig_loopback =8217;
7274: waveform_sig_loopback =3281;
7275: waveform_sig_loopback =6456;
7276: waveform_sig_loopback =8559;
7277: waveform_sig_loopback =5808;
7278: waveform_sig_loopback =5163;
7279: waveform_sig_loopback =5360;
7280: waveform_sig_loopback =7590;
7281: waveform_sig_loopback =6987;
7282: waveform_sig_loopback =4834;
7283: waveform_sig_loopback =6111;
7284: waveform_sig_loopback =6376;
7285: waveform_sig_loopback =6070;
7286: waveform_sig_loopback =6416;
7287: waveform_sig_loopback =4768;
7288: waveform_sig_loopback =7164;
7289: waveform_sig_loopback =5814;
7290: waveform_sig_loopback =5373;
7291: waveform_sig_loopback =6332;
7292: waveform_sig_loopback =5690;
7293: waveform_sig_loopback =5915;
7294: waveform_sig_loopback =5317;
7295: waveform_sig_loopback =6891;
7296: waveform_sig_loopback =4806;
7297: waveform_sig_loopback =5641;
7298: waveform_sig_loopback =6456;
7299: waveform_sig_loopback =5387;
7300: waveform_sig_loopback =4932;
7301: waveform_sig_loopback =6494;
7302: waveform_sig_loopback =5926;
7303: waveform_sig_loopback =4091;
7304: waveform_sig_loopback =6502;
7305: waveform_sig_loopback =6131;
7306: waveform_sig_loopback =4154;
7307: waveform_sig_loopback =5482;
7308: waveform_sig_loopback =6501;
7309: waveform_sig_loopback =5132;
7310: waveform_sig_loopback =4050;
7311: waveform_sig_loopback =6409;
7312: waveform_sig_loopback =5802;
7313: waveform_sig_loopback =4234;
7314: waveform_sig_loopback =7189;
7315: waveform_sig_loopback =2105;
7316: waveform_sig_loopback =5271;
7317: waveform_sig_loopback =7721;
7318: waveform_sig_loopback =4263;
7319: waveform_sig_loopback =4007;
7320: waveform_sig_loopback =4544;
7321: waveform_sig_loopback =6039;
7322: waveform_sig_loopback =6012;
7323: waveform_sig_loopback =3585;
7324: waveform_sig_loopback =4849;
7325: waveform_sig_loopback =5339;
7326: waveform_sig_loopback =4624;
7327: waveform_sig_loopback =5179;
7328: waveform_sig_loopback =3684;
7329: waveform_sig_loopback =5798;
7330: waveform_sig_loopback =4545;
7331: waveform_sig_loopback =4143;
7332: waveform_sig_loopback =4998;
7333: waveform_sig_loopback =4473;
7334: waveform_sig_loopback =4541;
7335: waveform_sig_loopback =3967;
7336: waveform_sig_loopback =5721;
7337: waveform_sig_loopback =3434;
7338: waveform_sig_loopback =4230;
7339: waveform_sig_loopback =5379;
7340: waveform_sig_loopback =3729;
7341: waveform_sig_loopback =3690;
7342: waveform_sig_loopback =5305;
7343: waveform_sig_loopback =3999;
7344: waveform_sig_loopback =3148;
7345: waveform_sig_loopback =4977;
7346: waveform_sig_loopback =4603;
7347: waveform_sig_loopback =2963;
7348: waveform_sig_loopback =3797;
7349: waveform_sig_loopback =5314;
7350: waveform_sig_loopback =3622;
7351: waveform_sig_loopback =2422;
7352: waveform_sig_loopback =5319;
7353: waveform_sig_loopback =3982;
7354: waveform_sig_loopback =2933;
7355: waveform_sig_loopback =5803;
7356: waveform_sig_loopback =235;
7357: waveform_sig_loopback =4166;
7358: waveform_sig_loopback =6153;
7359: waveform_sig_loopback =2601;
7360: waveform_sig_loopback =2592;
7361: waveform_sig_loopback =3076;
7362: waveform_sig_loopback =4483;
7363: waveform_sig_loopback =4561;
7364: waveform_sig_loopback =1770;
7365: waveform_sig_loopback =3400;
7366: waveform_sig_loopback =3905;
7367: waveform_sig_loopback =2908;
7368: waveform_sig_loopback =3702;
7369: waveform_sig_loopback =2165;
7370: waveform_sig_loopback =4108;
7371: waveform_sig_loopback =3039;
7372: waveform_sig_loopback =2563;
7373: waveform_sig_loopback =3286;
7374: waveform_sig_loopback =3164;
7375: waveform_sig_loopback =2666;
7376: waveform_sig_loopback =2501;
7377: waveform_sig_loopback =4221;
7378: waveform_sig_loopback =1424;
7379: waveform_sig_loopback =3017;
7380: waveform_sig_loopback =3546;
7381: waveform_sig_loopback =1976;
7382: waveform_sig_loopback =2356;
7383: waveform_sig_loopback =3394;
7384: waveform_sig_loopback =2445;
7385: waveform_sig_loopback =1563;
7386: waveform_sig_loopback =3215;
7387: waveform_sig_loopback =3035;
7388: waveform_sig_loopback =1231;
7389: waveform_sig_loopback =2160;
7390: waveform_sig_loopback =3761;
7391: waveform_sig_loopback =1713;
7392: waveform_sig_loopback =769;
7393: waveform_sig_loopback =3880;
7394: waveform_sig_loopback =1960;
7395: waveform_sig_loopback =1419;
7396: waveform_sig_loopback =4080;
7397: waveform_sig_loopback =-1756;
7398: waveform_sig_loopback =2963;
7399: waveform_sig_loopback =4153;
7400: waveform_sig_loopback =638;
7401: waveform_sig_loopback =1185;
7402: waveform_sig_loopback =1011;
7403: waveform_sig_loopback =2875;
7404: waveform_sig_loopback =2857;
7405: waveform_sig_loopback =-324;
7406: waveform_sig_loopback =2075;
7407: waveform_sig_loopback =1698;
7408: waveform_sig_loopback =1085;
7409: waveform_sig_loopback =2211;
7410: waveform_sig_loopback =92;
7411: waveform_sig_loopback =2366;
7412: waveform_sig_loopback =1084;
7413: waveform_sig_loopback =828;
7414: waveform_sig_loopback =1636;
7415: waveform_sig_loopback =1154;
7416: waveform_sig_loopback =619;
7417: waveform_sig_loopback =1085;
7418: waveform_sig_loopback =2245;
7419: waveform_sig_loopback =-627;
7420: waveform_sig_loopback =1412;
7421: waveform_sig_loopback =1472;
7422: waveform_sig_loopback =209;
7423: waveform_sig_loopback =541;
7424: waveform_sig_loopback =1326;
7425: waveform_sig_loopback =842;
7426: waveform_sig_loopback =-381;
7427: waveform_sig_loopback =1229;
7428: waveform_sig_loopback =1322;
7429: waveform_sig_loopback =-895;
7430: waveform_sig_loopback =426;
7431: waveform_sig_loopback =1914;
7432: waveform_sig_loopback =-555;
7433: waveform_sig_loopback =-726;
7434: waveform_sig_loopback =1934;
7435: waveform_sig_loopback =-310;
7436: waveform_sig_loopback =20;
7437: waveform_sig_loopback =1794;
7438: waveform_sig_loopback =-3681;
7439: waveform_sig_loopback =1450;
7440: waveform_sig_loopback =1817;
7441: waveform_sig_loopback =-1010;
7442: waveform_sig_loopback =-780;
7443: waveform_sig_loopback =-1043;
7444: waveform_sig_loopback =1435;
7445: waveform_sig_loopback =605;
7446: waveform_sig_loopback =-2236;
7447: waveform_sig_loopback =453;
7448: waveform_sig_loopback =-389;
7449: waveform_sig_loopback =-445;
7450: waveform_sig_loopback =56;
7451: waveform_sig_loopback =-1956;
7452: waveform_sig_loopback =951;
7453: waveform_sig_loopback =-997;
7454: waveform_sig_loopback =-1226;
7455: waveform_sig_loopback =-187;
7456: waveform_sig_loopback =-794;
7457: waveform_sig_loopback =-1139;
7458: waveform_sig_loopback =-840;
7459: waveform_sig_loopback =-1;
7460: waveform_sig_loopback =-2235;
7461: waveform_sig_loopback =-366;
7462: waveform_sig_loopback =-744;
7463: waveform_sig_loopback =-1461;
7464: waveform_sig_loopback =-1389;
7465: waveform_sig_loopback =-567;
7466: waveform_sig_loopback =-998;
7467: waveform_sig_loopback =-2572;
7468: waveform_sig_loopback =-273;
7469: waveform_sig_loopback =-658;
7470: waveform_sig_loopback =-3146;
7471: waveform_sig_loopback =-923;
7472: waveform_sig_loopback =-227;
7473: waveform_sig_loopback =-2470;
7474: waveform_sig_loopback =-2351;
7475: waveform_sig_loopback =-239;
7476: waveform_sig_loopback =-1939;
7477: waveform_sig_loopback =-1782;
7478: waveform_sig_loopback =-441;
7479: waveform_sig_loopback =-5290;
7480: waveform_sig_loopback =-406;
7481: waveform_sig_loopback =-170;
7482: waveform_sig_loopback =-2782;
7483: waveform_sig_loopback =-2920;
7484: waveform_sig_loopback =-2649;
7485: waveform_sig_loopback =-405;
7486: waveform_sig_loopback =-1573;
7487: waveform_sig_loopback =-3879;
7488: waveform_sig_loopback =-1403;
7489: waveform_sig_loopback =-2457;
7490: waveform_sig_loopback =-2030;
7491: waveform_sig_loopback =-2076;
7492: waveform_sig_loopback =-3716;
7493: waveform_sig_loopback =-726;
7494: waveform_sig_loopback =-3221;
7495: waveform_sig_loopback =-2778;
7496: waveform_sig_loopback =-2016;
7497: waveform_sig_loopback =-2880;
7498: waveform_sig_loopback =-2697;
7499: waveform_sig_loopback =-2770;
7500: waveform_sig_loopback =-1925;
7501: waveform_sig_loopback =-3795;
7502: waveform_sig_loopback =-2527;
7503: waveform_sig_loopback =-2317;
7504: waveform_sig_loopback =-3332;
7505: waveform_sig_loopback =-3432;
7506: waveform_sig_loopback =-1942;
7507: waveform_sig_loopback =-3218;
7508: waveform_sig_loopback =-4268;
7509: waveform_sig_loopback =-1860;
7510: waveform_sig_loopback =-2854;
7511: waveform_sig_loopback =-4693;
7512: waveform_sig_loopback =-2659;
7513: waveform_sig_loopback =-2208;
7514: waveform_sig_loopback =-4116;
7515: waveform_sig_loopback =-4204;
7516: waveform_sig_loopback =-2005;
7517: waveform_sig_loopback =-3717;
7518: waveform_sig_loopback =-3581;
7519: waveform_sig_loopback =-2278;
7520: waveform_sig_loopback =-6980;
7521: waveform_sig_loopback =-2130;
7522: waveform_sig_loopback =-1877;
7523: waveform_sig_loopback =-4537;
7524: waveform_sig_loopback =-4852;
7525: waveform_sig_loopback =-4014;
7526: waveform_sig_loopback =-2284;
7527: waveform_sig_loopback =-3454;
7528: waveform_sig_loopback =-5292;
7529: waveform_sig_loopback =-3422;
7530: waveform_sig_loopback =-3979;
7531: waveform_sig_loopback =-3721;
7532: waveform_sig_loopback =-4075;
7533: waveform_sig_loopback =-4919;
7534: waveform_sig_loopback =-2720;
7535: waveform_sig_loopback =-4900;
7536: waveform_sig_loopback =-4203;
7537: waveform_sig_loopback =-4036;
7538: waveform_sig_loopback =-4270;
7539: waveform_sig_loopback =-4461;
7540: waveform_sig_loopback =-4476;
7541: waveform_sig_loopback =-3385;
7542: waveform_sig_loopback =-5586;
7543: waveform_sig_loopback =-4107;
7544: waveform_sig_loopback =-3805;
7545: waveform_sig_loopback =-5132;
7546: waveform_sig_loopback =-4956;
7547: waveform_sig_loopback =-3427;
7548: waveform_sig_loopback =-5119;
7549: waveform_sig_loopback =-5588;
7550: waveform_sig_loopback =-3382;
7551: waveform_sig_loopback =-4693;
7552: waveform_sig_loopback =-5963;
7553: waveform_sig_loopback =-4319;
7554: waveform_sig_loopback =-3828;
7555: waveform_sig_loopback =-5516;
7556: waveform_sig_loopback =-6012;
7557: waveform_sig_loopback =-3203;
7558: waveform_sig_loopback =-5376;
7559: waveform_sig_loopback =-5177;
7560: waveform_sig_loopback =-3597;
7561: waveform_sig_loopback =-8718;
7562: waveform_sig_loopback =-3363;
7563: waveform_sig_loopback =-3349;
7564: waveform_sig_loopback =-6348;
7565: waveform_sig_loopback =-6048;
7566: waveform_sig_loopback =-5433;
7567: waveform_sig_loopback =-3926;
7568: waveform_sig_loopback =-4799;
7569: waveform_sig_loopback =-6802;
7570: waveform_sig_loopback =-4865;
7571: waveform_sig_loopback =-5182;
7572: waveform_sig_loopback =-5391;
7573: waveform_sig_loopback =-5398;
7574: waveform_sig_loopback =-6182;
7575: waveform_sig_loopback =-4430;
7576: waveform_sig_loopback =-6028;
7577: waveform_sig_loopback =-5667;
7578: waveform_sig_loopback =-5467;
7579: waveform_sig_loopback =-5416;
7580: waveform_sig_loopback =-6129;
7581: waveform_sig_loopback =-5610;
7582: waveform_sig_loopback =-4755;
7583: waveform_sig_loopback =-7180;
7584: waveform_sig_loopback =-5203;
7585: waveform_sig_loopback =-5168;
7586: waveform_sig_loopback =-6662;
7587: waveform_sig_loopback =-6012;
7588: waveform_sig_loopback =-4801;
7589: waveform_sig_loopback =-6551;
7590: waveform_sig_loopback =-6564;
7591: waveform_sig_loopback =-4943;
7592: waveform_sig_loopback =-5877;
7593: waveform_sig_loopback =-7084;
7594: waveform_sig_loopback =-5856;
7595: waveform_sig_loopback =-4674;
7596: waveform_sig_loopback =-7036;
7597: waveform_sig_loopback =-7206;
7598: waveform_sig_loopback =-4027;
7599: waveform_sig_loopback =-7163;
7600: waveform_sig_loopback =-5850;
7601: waveform_sig_loopback =-5061;
7602: waveform_sig_loopback =-10113;
7603: waveform_sig_loopback =-3905;
7604: waveform_sig_loopback =-5030;
7605: waveform_sig_loopback =-7468;
7606: waveform_sig_loopback =-6978;
7607: waveform_sig_loopback =-6814;
7608: waveform_sig_loopback =-4769;
7609: waveform_sig_loopback =-6057;
7610: waveform_sig_loopback =-8068;
7611: waveform_sig_loopback =-5677;
7612: waveform_sig_loopback =-6490;
7613: waveform_sig_loopback =-6370;
7614: waveform_sig_loopback =-6490;
7615: waveform_sig_loopback =-7302;
7616: waveform_sig_loopback =-5428;
7617: waveform_sig_loopback =-7039;
7618: waveform_sig_loopback =-6808;
7619: waveform_sig_loopback =-6490;
7620: waveform_sig_loopback =-6167;
7621: waveform_sig_loopback =-7477;
7622: waveform_sig_loopback =-6235;
7623: waveform_sig_loopback =-5859;
7624: waveform_sig_loopback =-8298;
7625: waveform_sig_loopback =-5580;
7626: waveform_sig_loopback =-6670;
7627: waveform_sig_loopback =-7301;
7628: waveform_sig_loopback =-6702;
7629: waveform_sig_loopback =-6122;
7630: waveform_sig_loopback =-7006;
7631: waveform_sig_loopback =-7699;
7632: waveform_sig_loopback =-5719;
7633: waveform_sig_loopback =-6553;
7634: waveform_sig_loopback =-8358;
7635: waveform_sig_loopback =-6237;
7636: waveform_sig_loopback =-5629;
7637: waveform_sig_loopback =-8102;
7638: waveform_sig_loopback =-7585;
7639: waveform_sig_loopback =-5015;
7640: waveform_sig_loopback =-8021;
7641: waveform_sig_loopback =-6276;
7642: waveform_sig_loopback =-6234;
7643: waveform_sig_loopback =-10641;
7644: waveform_sig_loopback =-4395;
7645: waveform_sig_loopback =-6047;
7646: waveform_sig_loopback =-7997;
7647: waveform_sig_loopback =-7743;
7648: waveform_sig_loopback =-7483;
7649: waveform_sig_loopback =-5225;
7650: waveform_sig_loopback =-6845;
7651: waveform_sig_loopback =-8812;
7652: waveform_sig_loopback =-5970;
7653: waveform_sig_loopback =-7400;
7654: waveform_sig_loopback =-6830;
7655: waveform_sig_loopback =-6957;
7656: waveform_sig_loopback =-8178;
7657: waveform_sig_loopback =-5597;
7658: waveform_sig_loopback =-7800;
7659: waveform_sig_loopback =-7468;
7660: waveform_sig_loopback =-6617;
7661: waveform_sig_loopback =-7181;
7662: waveform_sig_loopback =-7779;
7663: waveform_sig_loopback =-6492;
7664: waveform_sig_loopback =-6879;
7665: waveform_sig_loopback =-8236;
7666: waveform_sig_loopback =-6365;
7667: waveform_sig_loopback =-7129;
7668: waveform_sig_loopback =-7450;
7669: waveform_sig_loopback =-7606;
7670: waveform_sig_loopback =-6153;
7671: waveform_sig_loopback =-7604;
7672: waveform_sig_loopback =-8213;
7673: waveform_sig_loopback =-5835;
7674: waveform_sig_loopback =-7217;
7675: waveform_sig_loopback =-8580;
7676: waveform_sig_loopback =-6500;
7677: waveform_sig_loopback =-6136;
7678: waveform_sig_loopback =-8462;
7679: waveform_sig_loopback =-7779;
7680: waveform_sig_loopback =-5435;
7681: waveform_sig_loopback =-8419;
7682: waveform_sig_loopback =-6294;
7683: waveform_sig_loopback =-6912;
7684: waveform_sig_loopback =-10661;
7685: waveform_sig_loopback =-4532;
7686: waveform_sig_loopback =-6581;
7687: waveform_sig_loopback =-7917;
7688: waveform_sig_loopback =-8203;
7689: waveform_sig_loopback =-7605;
7690: waveform_sig_loopback =-5196;
7691: waveform_sig_loopback =-7508;
7692: waveform_sig_loopback =-8667;
7693: waveform_sig_loopback =-6154;
7694: waveform_sig_loopback =-7816;
7695: waveform_sig_loopback =-6508;
7696: waveform_sig_loopback =-7611;
7697: waveform_sig_loopback =-8032;
7698: waveform_sig_loopback =-5482;
7699: waveform_sig_loopback =-8361;
7700: waveform_sig_loopback =-7074;
7701: waveform_sig_loopback =-6930;
7702: waveform_sig_loopback =-7317;
7703: waveform_sig_loopback =-7436;
7704: waveform_sig_loopback =-6928;
7705: waveform_sig_loopback =-6695;
7706: waveform_sig_loopback =-8242;
7707: waveform_sig_loopback =-6497;
7708: waveform_sig_loopback =-6835;
7709: waveform_sig_loopback =-7725;
7710: waveform_sig_loopback =-7354;
7711: waveform_sig_loopback =-6067;
7712: waveform_sig_loopback =-7717;
7713: waveform_sig_loopback =-7941;
7714: waveform_sig_loopback =-5706;
7715: waveform_sig_loopback =-7221;
7716: waveform_sig_loopback =-8504;
7717: waveform_sig_loopback =-6146;
7718: waveform_sig_loopback =-6210;
7719: waveform_sig_loopback =-8282;
7720: waveform_sig_loopback =-7386;
7721: waveform_sig_loopback =-5512;
7722: waveform_sig_loopback =-8003;
7723: waveform_sig_loopback =-6007;
7724: waveform_sig_loopback =-7080;
7725: waveform_sig_loopback =-9939;
7726: waveform_sig_loopback =-4552;
7727: waveform_sig_loopback =-6219;
7728: waveform_sig_loopback =-7581;
7729: waveform_sig_loopback =-8336;
7730: waveform_sig_loopback =-6676;
7731: waveform_sig_loopback =-5251;
7732: waveform_sig_loopback =-7241;
7733: waveform_sig_loopback =-7972;
7734: waveform_sig_loopback =-6287;
7735: waveform_sig_loopback =-7011;
7736: waveform_sig_loopback =-6256;
7737: waveform_sig_loopback =-7476;
7738: waveform_sig_loopback =-7142;
7739: waveform_sig_loopback =-5555;
7740: waveform_sig_loopback =-7778;
7741: waveform_sig_loopback =-6512;
7742: waveform_sig_loopback =-6776;
7743: waveform_sig_loopback =-6501;
7744: waveform_sig_loopback =-7348;
7745: waveform_sig_loopback =-6199;
7746: waveform_sig_loopback =-6297;
7747: waveform_sig_loopback =-7813;
7748: waveform_sig_loopback =-5877;
7749: waveform_sig_loopback =-6443;
7750: waveform_sig_loopback =-7085;
7751: waveform_sig_loopback =-7009;
7752: waveform_sig_loopback =-5273;
7753: waveform_sig_loopback =-7473;
7754: waveform_sig_loopback =-7181;
7755: waveform_sig_loopback =-5126;
7756: waveform_sig_loopback =-7154;
7757: waveform_sig_loopback =-7244;
7758: waveform_sig_loopback =-5739;
7759: waveform_sig_loopback =-5798;
7760: waveform_sig_loopback =-7556;
7761: waveform_sig_loopback =-6817;
7762: waveform_sig_loopback =-4499;
7763: waveform_sig_loopback =-7655;
7764: waveform_sig_loopback =-5524;
7765: waveform_sig_loopback =-6053;
7766: waveform_sig_loopback =-9403;
7767: waveform_sig_loopback =-3778;
7768: waveform_sig_loopback =-5383;
7769: waveform_sig_loopback =-7268;
7770: waveform_sig_loopback =-7128;
7771: waveform_sig_loopback =-6090;
7772: waveform_sig_loopback =-4707;
7773: waveform_sig_loopback =-6095;
7774: waveform_sig_loopback =-7537;
7775: waveform_sig_loopback =-5300;
7776: waveform_sig_loopback =-6247;
7777: waveform_sig_loopback =-5593;
7778: waveform_sig_loopback =-6424;
7779: waveform_sig_loopback =-6394;
7780: waveform_sig_loopback =-4769;
7781: waveform_sig_loopback =-6783;
7782: waveform_sig_loopback =-5742;
7783: waveform_sig_loopback =-5890;
7784: waveform_sig_loopback =-5590;
7785: waveform_sig_loopback =-6446;
7786: waveform_sig_loopback =-5264;
7787: waveform_sig_loopback =-5387;
7788: waveform_sig_loopback =-6929;
7789: waveform_sig_loopback =-4862;
7790: waveform_sig_loopback =-5377;
7791: waveform_sig_loopback =-6478;
7792: waveform_sig_loopback =-5549;
7793: waveform_sig_loopback =-4519;
7794: waveform_sig_loopback =-6621;
7795: waveform_sig_loopback =-5797;
7796: waveform_sig_loopback =-4332;
7797: waveform_sig_loopback =-5846;
7798: waveform_sig_loopback =-6416;
7799: waveform_sig_loopback =-4789;
7800: waveform_sig_loopback =-4336;
7801: waveform_sig_loopback =-6658;
7802: waveform_sig_loopback =-5819;
7803: waveform_sig_loopback =-3276;
7804: waveform_sig_loopback =-6771;
7805: waveform_sig_loopback =-3940;
7806: waveform_sig_loopback =-5394;
7807: waveform_sig_loopback =-8392;
7808: waveform_sig_loopback =-2069;
7809: waveform_sig_loopback =-4674;
7810: waveform_sig_loopback =-6163;
7811: waveform_sig_loopback =-5776;
7812: waveform_sig_loopback =-5016;
7813: waveform_sig_loopback =-3276;
7814: waveform_sig_loopback =-5142;
7815: waveform_sig_loopback =-6385;
7816: waveform_sig_loopback =-3783;
7817: waveform_sig_loopback =-5237;
7818: waveform_sig_loopback =-4382;
7819: waveform_sig_loopback =-5127;
7820: waveform_sig_loopback =-5158;
7821: waveform_sig_loopback =-3494;
7822: waveform_sig_loopback =-5584;
7823: waveform_sig_loopback =-4445;
7824: waveform_sig_loopback =-4514;
7825: waveform_sig_loopback =-4291;
7826: waveform_sig_loopback =-5344;
7827: waveform_sig_loopback =-3710;
7828: waveform_sig_loopback =-4135;
7829: waveform_sig_loopback =-5789;
7830: waveform_sig_loopback =-3175;
7831: waveform_sig_loopback =-4365;
7832: waveform_sig_loopback =-5012;
7833: waveform_sig_loopback =-3922;
7834: waveform_sig_loopback =-3621;
7835: waveform_sig_loopback =-4814;
7836: waveform_sig_loopback =-4557;
7837: waveform_sig_loopback =-2991;
7838: waveform_sig_loopback =-4214;
7839: waveform_sig_loopback =-5404;
7840: waveform_sig_loopback =-2923;
7841: waveform_sig_loopback =-3086;
7842: waveform_sig_loopback =-5448;
7843: waveform_sig_loopback =-3921;
7844: waveform_sig_loopback =-2115;
7845: waveform_sig_loopback =-5279;
7846: waveform_sig_loopback =-2222;
7847: waveform_sig_loopback =-4246;
7848: waveform_sig_loopback =-6621;
7849: waveform_sig_loopback =-480;
7850: waveform_sig_loopback =-3409;
7851: waveform_sig_loopback =-4485;
7852: waveform_sig_loopback =-4303;
7853: waveform_sig_loopback =-3564;
7854: waveform_sig_loopback =-1545;
7855: waveform_sig_loopback =-3864;
7856: waveform_sig_loopback =-4810;
7857: waveform_sig_loopback =-2024;
7858: waveform_sig_loopback =-3959;
7859: waveform_sig_loopback =-2593;
7860: waveform_sig_loopback =-3673;
7861: waveform_sig_loopback =-3633;
7862: waveform_sig_loopback =-1684;
7863: waveform_sig_loopback =-4189;
7864: waveform_sig_loopback =-2823;
7865: waveform_sig_loopback =-2786;
7866: waveform_sig_loopback =-2900;
7867: waveform_sig_loopback =-3613;
7868: waveform_sig_loopback =-1973;
7869: waveform_sig_loopback =-2817;
7870: waveform_sig_loopback =-3823;
7871: waveform_sig_loopback =-1592;
7872: waveform_sig_loopback =-2897;
7873: waveform_sig_loopback =-3139;
7874: waveform_sig_loopback =-2397;
7875: waveform_sig_loopback =-1879;
7876: waveform_sig_loopback =-3096;
7877: waveform_sig_loopback =-3030;
7878: waveform_sig_loopback =-1093;
7879: waveform_sig_loopback =-2578;
7880: waveform_sig_loopback =-3836;
7881: waveform_sig_loopback =-852;
7882: waveform_sig_loopback =-1719;
7883: waveform_sig_loopback =-3680;
7884: waveform_sig_loopback =-1899;
7885: waveform_sig_loopback =-760;
7886: waveform_sig_loopback =-3313;
7887: waveform_sig_loopback =-445;
7888: waveform_sig_loopback =-2953;
7889: waveform_sig_loopback =-4399;
7890: waveform_sig_loopback =1127;
7891: waveform_sig_loopback =-1722;
7892: waveform_sig_loopback =-2572;
7893: waveform_sig_loopback =-2752;
7894: waveform_sig_loopback =-1528;
7895: waveform_sig_loopback =311;
7896: waveform_sig_loopback =-2413;
7897: waveform_sig_loopback =-2675;
7898: waveform_sig_loopback =-362;
7899: waveform_sig_loopback =-2224;
7900: waveform_sig_loopback =-541;
7901: waveform_sig_loopback =-2210;
7902: waveform_sig_loopback =-1578;
7903: waveform_sig_loopback =75;
7904: waveform_sig_loopback =-2558;
7905: waveform_sig_loopback =-793;
7906: waveform_sig_loopback =-1017;
7907: waveform_sig_loopback =-1184;
7908: waveform_sig_loopback =-1586;
7909: waveform_sig_loopback =-170;
7910: waveform_sig_loopback =-1203;
7911: waveform_sig_loopback =-1664;
7912: waveform_sig_loopback =-71;
7913: waveform_sig_loopback =-913;
7914: waveform_sig_loopback =-1198;
7915: waveform_sig_loopback =-856;
7916: waveform_sig_loopback =375;
7917: waveform_sig_loopback =-1614;
7918: waveform_sig_loopback =-1087;
7919: waveform_sig_loopback =1018;
7920: waveform_sig_loopback =-1263;
7921: waveform_sig_loopback =-1550;
7922: waveform_sig_loopback =915;
7923: waveform_sig_loopback =-77;
7924: waveform_sig_loopback =-1551;
7925: waveform_sig_loopback =-170;
7926: waveform_sig_loopback =1147;
7927: waveform_sig_loopback =-1442;
7928: waveform_sig_loopback =1451;
7929: waveform_sig_loopback =-1257;
7930: waveform_sig_loopback =-2297;
7931: waveform_sig_loopback =2943;
7932: waveform_sig_loopback =67;
7933: waveform_sig_loopback =-662;
7934: waveform_sig_loopback =-1043;
7935: waveform_sig_loopback =645;
7936: waveform_sig_loopback =2012;
7937: waveform_sig_loopback =-702;
7938: waveform_sig_loopback =-444;
7939: waveform_sig_loopback =1223;
7940: waveform_sig_loopback =-178;
7941: waveform_sig_loopback =1443;
7942: waveform_sig_loopback =-640;
7943: waveform_sig_loopback =735;
7944: waveform_sig_loopback =1723;
7945: waveform_sig_loopback =-698;
7946: waveform_sig_loopback =1358;
7947: waveform_sig_loopback =570;
7948: waveform_sig_loopback =851;
7949: waveform_sig_loopback =368;
7950: waveform_sig_loopback =1522;
7951: waveform_sig_loopback =887;
7952: waveform_sig_loopback =148;
7953: waveform_sig_loopback =1757;
7954: waveform_sig_loopback =1208;
7955: waveform_sig_loopback =380;
7956: waveform_sig_loopback =1279;
7957: waveform_sig_loopback =2212;
7958: waveform_sig_loopback =4;
7959: waveform_sig_loopback =1178;
7960: waveform_sig_loopback =2721;
7961: waveform_sig_loopback =509;
7962: waveform_sig_loopback =570;
7963: waveform_sig_loopback =2683;
7964: waveform_sig_loopback =1882;
7965: waveform_sig_loopback =292;
7966: waveform_sig_loopback =1725;
7967: waveform_sig_loopback =3045;
7968: waveform_sig_loopback =395;
7969: waveform_sig_loopback =3335;
7970: waveform_sig_loopback =443;
7971: waveform_sig_loopback =-233;
7972: waveform_sig_loopback =4767;
7973: waveform_sig_loopback =1965;
7974: waveform_sig_loopback =1046;
7975: waveform_sig_loopback =860;
7976: waveform_sig_loopback =2772;
7977: waveform_sig_loopback =3545;
7978: waveform_sig_loopback =1269;
7979: waveform_sig_loopback =1504;
7980: waveform_sig_loopback =2860;
7981: waveform_sig_loopback =2018;
7982: waveform_sig_loopback =2940;
7983: waveform_sig_loopback =1297;
7984: waveform_sig_loopback =2894;
7985: waveform_sig_loopback =3043;
7986: waveform_sig_loopback =1530;
7987: waveform_sig_loopback =3098;
7988: waveform_sig_loopback =2290;
7989: waveform_sig_loopback =2972;
7990: waveform_sig_loopback =1828;
7991: waveform_sig_loopback =3652;
7992: waveform_sig_loopback =2595;
7993: waveform_sig_loopback =1805;
7994: waveform_sig_loopback =3844;
7995: waveform_sig_loopback =2755;
7996: waveform_sig_loopback =2178;
7997: waveform_sig_loopback =3275;
7998: waveform_sig_loopback =3834;
7999: waveform_sig_loopback =1831;
8000: waveform_sig_loopback =3124;
8001: waveform_sig_loopback =4428;
8002: waveform_sig_loopback =2161;
8003: waveform_sig_loopback =2563;
8004: waveform_sig_loopback =4380;
8005: waveform_sig_loopback =3554;
8006: waveform_sig_loopback =2123;
8007: waveform_sig_loopback =3396;
8008: waveform_sig_loopback =5011;
8009: waveform_sig_loopback =1957;
8010: waveform_sig_loopback =5136;
8011: waveform_sig_loopback =2295;
8012: waveform_sig_loopback =1330;
8013: waveform_sig_loopback =6791;
8014: waveform_sig_loopback =3614;
8015: waveform_sig_loopback =2450;
8016: waveform_sig_loopback =3123;
8017: waveform_sig_loopback =4165;
8018: waveform_sig_loopback =5274;
8019: waveform_sig_loopback =3145;
8020: waveform_sig_loopback =2872;
8021: waveform_sig_loopback =4898;
8022: waveform_sig_loopback =3519;
8023: waveform_sig_loopback =4540;
8024: waveform_sig_loopback =3248;
8025: waveform_sig_loopback =4295;
8026: waveform_sig_loopback =4816;
8027: waveform_sig_loopback =3307;
8028: waveform_sig_loopback =4488;
8029: waveform_sig_loopback =4168;
8030: waveform_sig_loopback =4492;
8031: waveform_sig_loopback =3473;
8032: waveform_sig_loopback =5394;
8033: waveform_sig_loopback =4082;
8034: waveform_sig_loopback =3505;
8035: waveform_sig_loopback =5529;
8036: waveform_sig_loopback =4347;
8037: waveform_sig_loopback =3660;
8038: waveform_sig_loopback =5138;
8039: waveform_sig_loopback =5113;
8040: waveform_sig_loopback =3425;
8041: waveform_sig_loopback =4908;
8042: waveform_sig_loopback =5606;
8043: waveform_sig_loopback =4037;
8044: waveform_sig_loopback =3907;
8045: waveform_sig_loopback =5918;
8046: waveform_sig_loopback =5337;
8047: waveform_sig_loopback =3217;
8048: waveform_sig_loopback =5382;
8049: waveform_sig_loopback =6349;
8050: waveform_sig_loopback =3201;
8051: waveform_sig_loopback =7180;
8052: waveform_sig_loopback =3216;
8053: waveform_sig_loopback =3154;
8054: waveform_sig_loopback =8487;
8055: waveform_sig_loopback =4546;
8056: waveform_sig_loopback =4391;
8057: waveform_sig_loopback =4475;
8058: waveform_sig_loopback =5640;
8059: waveform_sig_loopback =7009;
8060: waveform_sig_loopback =4260;
8061: waveform_sig_loopback =4578;
8062: waveform_sig_loopback =6374;
8063: waveform_sig_loopback =4840;
8064: waveform_sig_loopback =6098;
8065: waveform_sig_loopback =4640;
8066: waveform_sig_loopback =5768;
8067: waveform_sig_loopback =6249;
8068: waveform_sig_loopback =4704;
8069: waveform_sig_loopback =5826;
8070: waveform_sig_loopback =5652;
8071: waveform_sig_loopback =5742;
8072: waveform_sig_loopback =4755;
8073: waveform_sig_loopback =7010;
8074: waveform_sig_loopback =4992;
8075: waveform_sig_loopback =5034;
8076: waveform_sig_loopback =6936;
8077: waveform_sig_loopback =5235;
8078: waveform_sig_loopback =5376;
8079: waveform_sig_loopback =6267;
8080: waveform_sig_loopback =6281;
8081: waveform_sig_loopback =5023;
8082: waveform_sig_loopback =5887;
8083: waveform_sig_loopback =7038;
8084: waveform_sig_loopback =5243;
8085: waveform_sig_loopback =5020;
8086: waveform_sig_loopback =7535;
8087: waveform_sig_loopback =6264;
8088: waveform_sig_loopback =4423;
8089: waveform_sig_loopback =7008;
8090: waveform_sig_loopback =7130;
8091: waveform_sig_loopback =4693;
8092: waveform_sig_loopback =8465;
8093: waveform_sig_loopback =3846;
8094: waveform_sig_loopback =4989;
8095: waveform_sig_loopback =9361;
8096: waveform_sig_loopback =5685;
8097: waveform_sig_loopback =5657;
8098: waveform_sig_loopback =5268;
8099: waveform_sig_loopback =6999;
8100: waveform_sig_loopback =8075;
8101: waveform_sig_loopback =5128;
8102: waveform_sig_loopback =5771;
8103: waveform_sig_loopback =7205;
8104: waveform_sig_loopback =5936;
8105: waveform_sig_loopback =7319;
8106: waveform_sig_loopback =5369;
8107: waveform_sig_loopback =6573;
8108: waveform_sig_loopback =7534;
8109: waveform_sig_loopback =5582;
8110: waveform_sig_loopback =6746;
8111: waveform_sig_loopback =6677;
8112: waveform_sig_loopback =6389;
8113: waveform_sig_loopback =6230;
8114: waveform_sig_loopback =7762;
8115: waveform_sig_loopback =5572;
8116: waveform_sig_loopback =6630;
8117: waveform_sig_loopback =7399;
8118: waveform_sig_loopback =6393;
8119: waveform_sig_loopback =6254;
8120: waveform_sig_loopback =6896;
8121: waveform_sig_loopback =7725;
8122: waveform_sig_loopback =5369;
8123: waveform_sig_loopback =7003;
8124: waveform_sig_loopback =8126;
8125: waveform_sig_loopback =5728;
8126: waveform_sig_loopback =6184;
8127: waveform_sig_loopback =8149;
8128: waveform_sig_loopback =7060;
8129: waveform_sig_loopback =5264;
8130: waveform_sig_loopback =7777;
8131: waveform_sig_loopback =7751;
8132: waveform_sig_loopback =5564;
8133: waveform_sig_loopback =9277;
8134: waveform_sig_loopback =4126;
8135: waveform_sig_loopback =6203;
8136: waveform_sig_loopback =9833;
8137: waveform_sig_loopback =6238;
8138: waveform_sig_loopback =6506;
8139: waveform_sig_loopback =5710;
8140: waveform_sig_loopback =8048;
8141: waveform_sig_loopback =8522;
8142: waveform_sig_loopback =5445;
8143: waveform_sig_loopback =6982;
8144: waveform_sig_loopback =7632;
8145: waveform_sig_loopback =6545;
8146: waveform_sig_loopback =7984;
8147: waveform_sig_loopback =5674;
8148: waveform_sig_loopback =7874;
8149: waveform_sig_loopback =7674;
8150: waveform_sig_loopback =5906;
8151: waveform_sig_loopback =7852;
8152: waveform_sig_loopback =6983;
8153: waveform_sig_loopback =7091;
8154: waveform_sig_loopback =6716;
8155: waveform_sig_loopback =8094;
8156: waveform_sig_loopback =6498;
8157: waveform_sig_loopback =6872;
8158: waveform_sig_loopback =7830;
8159: waveform_sig_loopback =7033;
8160: waveform_sig_loopback =6582;
8161: waveform_sig_loopback =7583;
8162: waveform_sig_loopback =7947;
8163: waveform_sig_loopback =5759;
8164: waveform_sig_loopback =7605;
8165: waveform_sig_loopback =8336;
8166: waveform_sig_loopback =5929;
8167: waveform_sig_loopback =6755;
8168: waveform_sig_loopback =8553;
8169: waveform_sig_loopback =7065;
8170: waveform_sig_loopback =5814;
8171: waveform_sig_loopback =8097;
8172: waveform_sig_loopback =7922;
8173: waveform_sig_loopback =6126;
8174: waveform_sig_loopback =9218;
8175: waveform_sig_loopback =4530;
8176: waveform_sig_loopback =6705;
8177: waveform_sig_loopback =9736;
8178: waveform_sig_loopback =6860;
8179: waveform_sig_loopback =6359;
8180: waveform_sig_loopback =6069;
8181: waveform_sig_loopback =8557;
8182: waveform_sig_loopback =8222;
8183: waveform_sig_loopback =6017;
8184: waveform_sig_loopback =7045;
8185: waveform_sig_loopback =7598;
8186: waveform_sig_loopback =7107;
8187: waveform_sig_loopback =7746;
8188: waveform_sig_loopback =5945;
8189: waveform_sig_loopback =8211;
8190: waveform_sig_loopback =7335;
8191: waveform_sig_loopback =6430;
8192: waveform_sig_loopback =7701;
8193: waveform_sig_loopback =6976;
8194: waveform_sig_loopback =7345;
8195: waveform_sig_loopback =6475;
8196: waveform_sig_loopback =8377;
8197: waveform_sig_loopback =6420;
8198: waveform_sig_loopback =6809;
8199: waveform_sig_loopback =7965;
8200: waveform_sig_loopback =6943;
8201: waveform_sig_loopback =6522;
8202: waveform_sig_loopback =7678;
8203: waveform_sig_loopback =7766;
8204: waveform_sig_loopback =5566;
8205: waveform_sig_loopback =7816;
8206: waveform_sig_loopback =8111;
8207: waveform_sig_loopback =5749;
8208: waveform_sig_loopback =6865;
8209: waveform_sig_loopback =8138;
8210: waveform_sig_loopback =7077;
8211: waveform_sig_loopback =5764;
8212: waveform_sig_loopback =7716;
8213: waveform_sig_loopback =8016;
8214: waveform_sig_loopback =5716;
8215: waveform_sig_loopback =9075;
8216: waveform_sig_loopback =4469;
8217: waveform_sig_loopback =6229;
8218: waveform_sig_loopback =9937;
8219: waveform_sig_loopback =6386;
8220: waveform_sig_loopback =5844;
8221: waveform_sig_loopback =6369;
8222: waveform_sig_loopback =7715;
8223: waveform_sig_loopback =8140;
8224: waveform_sig_loopback =5738;
8225: waveform_sig_loopback =6433;
8226: waveform_sig_loopback =7654;
8227: waveform_sig_loopback =6513;
8228: waveform_sig_loopback =7381;
8229: waveform_sig_loopback =5813;
8230: waveform_sig_loopback =7592;
8231: waveform_sig_loopback =7083;
8232: waveform_sig_loopback =6026;
8233: waveform_sig_loopback =7216;
8234: waveform_sig_loopback =6706;
8235: waveform_sig_loopback =6790;
8236: waveform_sig_loopback =6106;
8237: waveform_sig_loopback =7872;
8238: waveform_sig_loopback =5914;
8239: waveform_sig_loopback =6227;
8240: waveform_sig_loopback =7701;
8241: waveform_sig_loopback =6302;
8242: waveform_sig_loopback =5864;
8243: waveform_sig_loopback =7574;
8244: waveform_sig_loopback =6704;
8245: waveform_sig_loopback =5426;
8246: waveform_sig_loopback =7257;
8247: waveform_sig_loopback =7142;
8248: waveform_sig_loopback =5565;
8249: waveform_sig_loopback =5982;
8250: waveform_sig_loopback =7757;
8251: waveform_sig_loopback =6425;
8252: waveform_sig_loopback =4751;
8253: waveform_sig_loopback =7600;
8254: waveform_sig_loopback =7047;
8255: waveform_sig_loopback =5034;
8256: waveform_sig_loopback =8677;
8257: waveform_sig_loopback =3246;
8258: waveform_sig_loopback =5963;
8259: waveform_sig_loopback =9174;
8260: waveform_sig_loopback =5295;
8261: waveform_sig_loopback =5391;
8262: waveform_sig_loopback =5543;
8263: waveform_sig_loopback =7022;
8264: waveform_sig_loopback =7546;
8265: waveform_sig_loopback =4645;
8266: waveform_sig_loopback =5863;
8267: waveform_sig_loopback =6847;
8268: waveform_sig_loopback =5545;
8269: waveform_sig_loopback =6657;
8270: waveform_sig_loopback =4946;
8271: waveform_sig_loopback =6753;
8272: waveform_sig_loopback =6215;
8273: waveform_sig_loopback =5182;
8274: waveform_sig_loopback =6207;
8275: waveform_sig_loopback =5981;
8276: waveform_sig_loopback =5768;
8277: waveform_sig_loopback =5181;
8278: waveform_sig_loopback =7183;
8279: waveform_sig_loopback =4568;
8280: waveform_sig_loopback =5643;
8281: waveform_sig_loopback =6701;
8282: waveform_sig_loopback =4979;
8283: waveform_sig_loopback =5297;
8284: waveform_sig_loopback =6340;
8285: waveform_sig_loopback =5696;
8286: waveform_sig_loopback =4579;
8287: waveform_sig_loopback =5996;
8288: waveform_sig_loopback =6385;
8289: waveform_sig_loopback =4417;
8290: waveform_sig_loopback =4903;
8291: waveform_sig_loopback =6986;
8292: waveform_sig_loopback =5052;
8293: waveform_sig_loopback =3757;
8294: waveform_sig_loopback =6765;
8295: waveform_sig_loopback =5497;
8296: waveform_sig_loopback =4236;
8297: waveform_sig_loopback =7452;
8298: waveform_sig_loopback =1799;
8299: waveform_sig_loopback =5401;
8300: waveform_sig_loopback =7705;
8301: waveform_sig_loopback =4116;
8302: waveform_sig_loopback =4393;
8303: waveform_sig_loopback =4111;
8304: waveform_sig_loopback =6072;
8305: waveform_sig_loopback =6303;
8306: waveform_sig_loopback =3209;
8307: waveform_sig_loopback =4950;
8308: waveform_sig_loopback =5446;
8309: waveform_sig_loopback =4367;
8310: waveform_sig_loopback =5506;
8311: waveform_sig_loopback =3500;
8312: waveform_sig_loopback =5683;
8313: waveform_sig_loopback =4915;
8314: waveform_sig_loopback =3763;
8315: waveform_sig_loopback =5096;
8316: waveform_sig_loopback =4704;
8317: waveform_sig_loopback =4206;
8318: waveform_sig_loopback =4140;
8319: waveform_sig_loopback =5755;
8320: waveform_sig_loopback =3130;
8321: waveform_sig_loopback =4617;
8322: waveform_sig_loopback =5023;
8323: waveform_sig_loopback =3802;
8324: waveform_sig_loopback =3997;
8325: waveform_sig_loopback =4706;
8326: waveform_sig_loopback =4626;
8327: waveform_sig_loopback =2973;
8328: waveform_sig_loopback =4645;
8329: waveform_sig_loopback =5167;
8330: waveform_sig_loopback =2611;
8331: waveform_sig_loopback =3795;
8332: waveform_sig_loopback =5535;
8333: waveform_sig_loopback =3346;
8334: waveform_sig_loopback =2634;
8335: waveform_sig_loopback =5213;
8336: waveform_sig_loopback =3932;
8337: waveform_sig_loopback =3064;
8338: waveform_sig_loopback =5701;
8339: waveform_sig_loopback =286;
8340: waveform_sig_loopback =4233;
8341: waveform_sig_loopback =5938;
8342: waveform_sig_loopback =2726;
8343: waveform_sig_loopback =2857;
8344: waveform_sig_loopback =2520;
8345: waveform_sig_loopback =4843;
8346: waveform_sig_loopback =4529;
8347: waveform_sig_loopback =1598;
8348: waveform_sig_loopback =3732;
8349: waveform_sig_loopback =3561;
8350: waveform_sig_loopback =3037;
8351: waveform_sig_loopback =3867;
8352: waveform_sig_loopback =1721;
8353: waveform_sig_loopback =4413;
8354: waveform_sig_loopback =3028;
8355: waveform_sig_loopback =2211;
8356: waveform_sig_loopback =3599;
8357: waveform_sig_loopback =2876;
8358: waveform_sig_loopback =2653;
8359: waveform_sig_loopback =2651;
8360: waveform_sig_loopback =3825;
8361: waveform_sig_loopback =1650;
8362: waveform_sig_loopback =3030;
8363: waveform_sig_loopback =3159;
8364: waveform_sig_loopback =2373;
8365: waveform_sig_loopback =2128;
8366: waveform_sig_loopback =3172;
8367: waveform_sig_loopback =2936;
8368: waveform_sig_loopback =1007;
8369: waveform_sig_loopback =3306;
8370: waveform_sig_loopback =3294;
8371: waveform_sig_loopback =742;
8372: waveform_sig_loopback =2489;
8373: waveform_sig_loopback =3558;
8374: waveform_sig_loopback =1613;
8375: waveform_sig_loopback =1117;
8376: waveform_sig_loopback =3327;
8377: waveform_sig_loopback =2349;
8378: waveform_sig_loopback =1352;
8379: waveform_sig_loopback =3829;
8380: waveform_sig_loopback =-1328;
8381: waveform_sig_loopback =2520;
8382: waveform_sig_loopback =4181;
8383: waveform_sig_loopback =953;
8384: waveform_sig_loopback =984;
8385: waveform_sig_loopback =925;
8386: waveform_sig_loopback =3055;
8387: waveform_sig_loopback =2598;
8388: waveform_sig_loopback =-135;
8389: waveform_sig_loopback =2034;
8390: waveform_sig_loopback =1555;
8391: waveform_sig_loopback =1463;
8392: waveform_sig_loopback =1941;
8393: waveform_sig_loopback =-120;
8394: waveform_sig_loopback =2866;
8395: waveform_sig_loopback =847;
8396: waveform_sig_loopback =749;
8397: waveform_sig_loopback =1758;
8398: waveform_sig_loopback =808;
8399: waveform_sig_loopback =1149;
8400: waveform_sig_loopback =765;
8401: waveform_sig_loopback =1982;
8402: waveform_sig_loopback =12;
8403: waveform_sig_loopback =842;
8404: waveform_sig_loopback =1723;
8405: waveform_sig_loopback =421;
8406: waveform_sig_loopback =101;
8407: waveform_sig_loopback =1794;
8408: waveform_sig_loopback =662;
8409: waveform_sig_loopback =-528;
8410: waveform_sig_loopback =1549;
8411: waveform_sig_loopback =1184;
8412: waveform_sig_loopback =-858;
8413: waveform_sig_loopback =576;
8414: waveform_sig_loopback =1741;
8415: waveform_sig_loopback =-230;
8416: waveform_sig_loopback =-734;
8417: waveform_sig_loopback =1532;
8418: waveform_sig_loopback =380;
8419: waveform_sig_loopback =-379;
8420: waveform_sig_loopback =1823;
8421: waveform_sig_loopback =-3172;
8422: waveform_sig_loopback =766;
8423: waveform_sig_loopback =2255;
8424: waveform_sig_loopback =-928;
8425: waveform_sig_loopback =-1088;
8426: waveform_sig_loopback =-621;
8427: waveform_sig_loopback =1121;
8428: waveform_sig_loopback =538;
8429: waveform_sig_loopback =-1744;
8430: waveform_sig_loopback =-17;
8431: waveform_sig_loopback =-236;
8432: waveform_sig_loopback =-284;
8433: waveform_sig_loopback =-277;
8434: waveform_sig_loopback =-1520;
8435: waveform_sig_loopback =762;
8436: waveform_sig_loopback =-1149;
8437: waveform_sig_loopback =-773;
8438: waveform_sig_loopback =-464;
8439: waveform_sig_loopback =-731;
8440: waveform_sig_loopback =-874;
8441: waveform_sig_loopback =-1310;
8442: waveform_sig_loopback =488;
8443: waveform_sig_loopback =-2255;
8444: waveform_sig_loopback =-799;
8445: waveform_sig_loopback =-151;
8446: waveform_sig_loopback =-1720;
8447: waveform_sig_loopback =-1500;
8448: waveform_sig_loopback =-215;
8449: waveform_sig_loopback =-1320;
8450: waveform_sig_loopback =-2265;
8451: waveform_sig_loopback =-520;
8452: waveform_sig_loopback =-796;
8453: waveform_sig_loopback =-2583;
8454: waveform_sig_loopback =-1270;
8455: waveform_sig_loopback =-434;
8456: waveform_sig_loopback =-2136;
8457: waveform_sig_loopback =-2501;
8458: waveform_sig_loopback =-230;
8459: waveform_sig_loopback =-1704;
8460: waveform_sig_loopback =-2387;
8461: waveform_sig_loopback =199;
8462: waveform_sig_loopback =-5257;
8463: waveform_sig_loopback =-1076;
8464: waveform_sig_loopback =454;
8465: waveform_sig_loopback =-3040;
8466: waveform_sig_loopback =-2866;
8467: waveform_sig_loopback =-2448;
8468: waveform_sig_loopback =-958;
8469: waveform_sig_loopback =-1035;
8470: waveform_sig_loopback =-3836;
8471: waveform_sig_loopback =-2000;
8472: waveform_sig_loopback =-1774;
8473: waveform_sig_loopback =-2434;
8474: waveform_sig_loopback =-2031;
8475: waveform_sig_loopback =-3387;
8476: waveform_sig_loopback =-1334;
8477: waveform_sig_loopback =-2606;
8478: waveform_sig_loopback =-2991;
8479: waveform_sig_loopback =-2347;
8480: waveform_sig_loopback =-2334;
8481: waveform_sig_loopback =-3079;
8482: waveform_sig_loopback =-2772;
8483: waveform_sig_loopback =-1654;
8484: waveform_sig_loopback =-4112;
8485: waveform_sig_loopback =-2368;
8486: waveform_sig_loopback =-2264;
8487: waveform_sig_loopback =-3480;
8488: waveform_sig_loopback =-3295;
8489: waveform_sig_loopback =-1979;
8490: waveform_sig_loopback =-3306;
8491: waveform_sig_loopback =-4021;
8492: waveform_sig_loopback =-2055;
8493: waveform_sig_loopback =-2842;
8494: waveform_sig_loopback =-4359;
8495: waveform_sig_loopback =-3196;
8496: waveform_sig_loopback =-1919;
8497: waveform_sig_loopback =-3888;
8498: waveform_sig_loopback =-4815;
8499: waveform_sig_loopback =-1418;
8500: waveform_sig_loopback =-3954;
8501: waveform_sig_loopback =-3751;
8502: waveform_sig_loopback =-1709;
8503: waveform_sig_loopback =-7578;
8504: waveform_sig_loopback =-1790;
8505: waveform_sig_loopback =-1815;
8506: waveform_sig_loopback =-4929;
8507: waveform_sig_loopback =-4245;
8508: waveform_sig_loopback =-4433;
8509: waveform_sig_loopback =-2318;
8510: waveform_sig_loopback =-3059;
8511: waveform_sig_loopback =-5708;
8512: waveform_sig_loopback =-3198;
8513: waveform_sig_loopback =-3890;
8514: waveform_sig_loopback =-4106;
8515: waveform_sig_loopback =-3551;
8516: waveform_sig_loopback =-5212;
8517: waveform_sig_loopback =-2880;
8518: waveform_sig_loopback =-4478;
8519: waveform_sig_loopback =-4518;
8520: waveform_sig_loopback =-3902;
8521: waveform_sig_loopback =-4142;
8522: waveform_sig_loopback =-4769;
8523: waveform_sig_loopback =-4248;
8524: waveform_sig_loopback =-3267;
8525: waveform_sig_loopback =-5958;
8526: waveform_sig_loopback =-3730;
8527: waveform_sig_loopback =-3967;
8528: waveform_sig_loopback =-5169;
8529: waveform_sig_loopback =-4619;
8530: waveform_sig_loopback =-3899;
8531: waveform_sig_loopback =-4815;
8532: waveform_sig_loopback =-5515;
8533: waveform_sig_loopback =-3819;
8534: waveform_sig_loopback =-4182;
8535: waveform_sig_loopback =-6180;
8536: waveform_sig_loopback =-4595;
8537: waveform_sig_loopback =-3292;
8538: waveform_sig_loopback =-5954;
8539: waveform_sig_loopback =-5935;
8540: waveform_sig_loopback =-2953;
8541: waveform_sig_loopback =-5813;
8542: waveform_sig_loopback =-4863;
8543: waveform_sig_loopback =-3573;
8544: waveform_sig_loopback =-8903;
8545: waveform_sig_loopback =-3198;
8546: waveform_sig_loopback =-3669;
8547: waveform_sig_loopback =-6015;
8548: waveform_sig_loopback =-5938;
8549: waveform_sig_loopback =-5963;
8550: waveform_sig_loopback =-3492;
8551: waveform_sig_loopback =-4707;
8552: waveform_sig_loopback =-7183;
8553: waveform_sig_loopback =-4567;
8554: waveform_sig_loopback =-5313;
8555: waveform_sig_loopback =-5405;
8556: waveform_sig_loopback =-5159;
8557: waveform_sig_loopback =-6606;
8558: waveform_sig_loopback =-4096;
8559: waveform_sig_loopback =-5914;
8560: waveform_sig_loopback =-6085;
8561: waveform_sig_loopback =-5124;
8562: waveform_sig_loopback =-5452;
8563: waveform_sig_loopback =-6300;
8564: waveform_sig_loopback =-5271;
8565: waveform_sig_loopback =-5043;
8566: waveform_sig_loopback =-7098;
8567: waveform_sig_loopback =-4896;
8568: waveform_sig_loopback =-5743;
8569: waveform_sig_loopback =-6144;
8570: waveform_sig_loopback =-6167;
8571: waveform_sig_loopback =-5053;
8572: waveform_sig_loopback =-5926;
8573: waveform_sig_loopback =-7212;
8574: waveform_sig_loopback =-4650;
8575: waveform_sig_loopback =-5580;
8576: waveform_sig_loopback =-7638;
8577: waveform_sig_loopback =-5480;
8578: waveform_sig_loopback =-4754;
8579: waveform_sig_loopback =-7183;
8580: waveform_sig_loopback =-6977;
8581: waveform_sig_loopback =-4344;
8582: waveform_sig_loopback =-6936;
8583: waveform_sig_loopback =-5909;
8584: waveform_sig_loopback =-5164;
8585: waveform_sig_loopback =-9829;
8586: waveform_sig_loopback =-4139;
8587: waveform_sig_loopback =-5104;
8588: waveform_sig_loopback =-7090;
8589: waveform_sig_loopback =-7165;
8590: waveform_sig_loopback =-7011;
8591: waveform_sig_loopback =-4477;
8592: waveform_sig_loopback =-6130;
8593: waveform_sig_loopback =-8128;
8594: waveform_sig_loopback =-5425;
8595: waveform_sig_loopback =-6803;
8596: waveform_sig_loopback =-6091;
8597: waveform_sig_loopback =-6375;
8598: waveform_sig_loopback =-7697;
8599: waveform_sig_loopback =-4778;
8600: waveform_sig_loopback =-7423;
8601: waveform_sig_loopback =-6771;
8602: waveform_sig_loopback =-6056;
8603: waveform_sig_loopback =-6891;
8604: waveform_sig_loopback =-6849;
8605: waveform_sig_loopback =-6435;
8606: waveform_sig_loopback =-6104;
8607: waveform_sig_loopback =-7770;
8608: waveform_sig_loopback =-6154;
8609: waveform_sig_loopback =-6382;
8610: waveform_sig_loopback =-7201;
8611: waveform_sig_loopback =-7212;
8612: waveform_sig_loopback =-5652;
8613: waveform_sig_loopback =-7123;
8614: waveform_sig_loopback =-7995;
8615: waveform_sig_loopback =-5407;
8616: waveform_sig_loopback =-6655;
8617: waveform_sig_loopback =-8424;
8618: waveform_sig_loopback =-6178;
8619: waveform_sig_loopback =-5746;
8620: waveform_sig_loopback =-7986;
8621: waveform_sig_loopback =-7563;
8622: waveform_sig_loopback =-5320;
8623: waveform_sig_loopback =-7597;
8624: waveform_sig_loopback =-6495;
8625: waveform_sig_loopback =-6293;
8626: waveform_sig_loopback =-10203;
8627: waveform_sig_loopback =-4951;
8628: waveform_sig_loopback =-5848;
8629: waveform_sig_loopback =-7579;
8630: waveform_sig_loopback =-8278;
8631: waveform_sig_loopback =-7193;
8632: waveform_sig_loopback =-5254;
8633: waveform_sig_loopback =-7091;
8634: waveform_sig_loopback =-8344;
8635: waveform_sig_loopback =-6460;
8636: waveform_sig_loopback =-7188;
8637: waveform_sig_loopback =-6635;
8638: waveform_sig_loopback =-7421;
8639: waveform_sig_loopback =-7785;
8640: waveform_sig_loopback =-5660;
8641: waveform_sig_loopback =-8074;
8642: waveform_sig_loopback =-7034;
8643: waveform_sig_loopback =-6905;
8644: waveform_sig_loopback =-7176;
8645: waveform_sig_loopback =-7475;
8646: waveform_sig_loopback =-6948;
8647: waveform_sig_loopback =-6537;
8648: waveform_sig_loopback =-8302;
8649: waveform_sig_loopback =-6612;
8650: waveform_sig_loopback =-6749;
8651: waveform_sig_loopback =-7696;
8652: waveform_sig_loopback =-7665;
8653: waveform_sig_loopback =-5897;
8654: waveform_sig_loopback =-7841;
8655: waveform_sig_loopback =-8201;
8656: waveform_sig_loopback =-5639;
8657: waveform_sig_loopback =-7435;
8658: waveform_sig_loopback =-8462;
8659: waveform_sig_loopback =-6526;
8660: waveform_sig_loopback =-6303;
8661: waveform_sig_loopback =-8090;
8662: waveform_sig_loopback =-8128;
8663: waveform_sig_loopback =-5449;
8664: waveform_sig_loopback =-7932;
8665: waveform_sig_loopback =-6937;
8666: waveform_sig_loopback =-6380;
8667: waveform_sig_loopback =-10604;
8668: waveform_sig_loopback =-5172;
8669: waveform_sig_loopback =-5901;
8670: waveform_sig_loopback =-8208;
8671: waveform_sig_loopback =-8305;
8672: waveform_sig_loopback =-7224;
8673: waveform_sig_loopback =-5771;
8674: waveform_sig_loopback =-6989;
8675: waveform_sig_loopback =-8682;
8676: waveform_sig_loopback =-6637;
8677: waveform_sig_loopback =-7150;
8678: waveform_sig_loopback =-7009;
8679: waveform_sig_loopback =-7424;
8680: waveform_sig_loopback =-7783;
8681: waveform_sig_loopback =-5989;
8682: waveform_sig_loopback =-7951;
8683: waveform_sig_loopback =-7149;
8684: waveform_sig_loopback =-7045;
8685: waveform_sig_loopback =-7069;
8686: waveform_sig_loopback =-7592;
8687: waveform_sig_loopback =-6926;
8688: waveform_sig_loopback =-6547;
8689: waveform_sig_loopback =-8374;
8690: waveform_sig_loopback =-6600;
8691: waveform_sig_loopback =-6586;
8692: waveform_sig_loopback =-8003;
8693: waveform_sig_loopback =-7304;
8694: waveform_sig_loopback =-5846;
8695: waveform_sig_loopback =-8169;
8696: waveform_sig_loopback =-7588;
8697: waveform_sig_loopback =-5896;
8698: waveform_sig_loopback =-7325;
8699: waveform_sig_loopback =-8156;
8700: waveform_sig_loopback =-6718;
8701: waveform_sig_loopback =-5812;
8702: waveform_sig_loopback =-8173;
8703: waveform_sig_loopback =-7975;
8704: waveform_sig_loopback =-4953;
8705: waveform_sig_loopback =-8194;
8706: waveform_sig_loopback =-6410;
8707: waveform_sig_loopback =-6358;
8708: waveform_sig_loopback =-10595;
8709: waveform_sig_loopback =-4433;
8710: waveform_sig_loopback =-5977;
8711: waveform_sig_loopback =-8074;
8712: waveform_sig_loopback =-7756;
8713: waveform_sig_loopback =-7109;
8714: waveform_sig_loopback =-5362;
8715: waveform_sig_loopback =-6737;
8716: waveform_sig_loopback =-8536;
8717: waveform_sig_loopback =-6029;
8718: waveform_sig_loopback =-6921;
8719: waveform_sig_loopback =-6675;
8720: waveform_sig_loopback =-7027;
8721: waveform_sig_loopback =-7408;
8722: waveform_sig_loopback =-5653;
8723: waveform_sig_loopback =-7507;
8724: waveform_sig_loopback =-6766;
8725: waveform_sig_loopback =-6703;
8726: waveform_sig_loopback =-6476;
8727: waveform_sig_loopback =-7496;
8728: waveform_sig_loopback =-6218;
8729: waveform_sig_loopback =-6046;
8730: waveform_sig_loopback =-8229;
8731: waveform_sig_loopback =-5611;
8732: waveform_sig_loopback =-6454;
8733: waveform_sig_loopback =-7439;
8734: waveform_sig_loopback =-6422;
8735: waveform_sig_loopback =-5830;
8736: waveform_sig_loopback =-7211;
8737: waveform_sig_loopback =-7132;
8738: waveform_sig_loopback =-5462;
8739: waveform_sig_loopback =-6432;
8740: waveform_sig_loopback =-7921;
8741: waveform_sig_loopback =-5767;
8742: waveform_sig_loopback =-5242;
8743: waveform_sig_loopback =-7841;
8744: waveform_sig_loopback =-6887;
8745: waveform_sig_loopback =-4414;
8746: waveform_sig_loopback =-7702;
8747: waveform_sig_loopback =-5408;
8748: waveform_sig_loopback =-6007;
8749: waveform_sig_loopback =-9664;
8750: waveform_sig_loopback =-3542;
8751: waveform_sig_loopback =-5531;
8752: waveform_sig_loopback =-7229;
8753: waveform_sig_loopback =-6870;
8754: waveform_sig_loopback =-6544;
8755: waveform_sig_loopback =-4313;
8756: waveform_sig_loopback =-6093;
8757: waveform_sig_loopback =-7848;
8758: waveform_sig_loopback =-4853;
8759: waveform_sig_loopback =-6472;
8760: waveform_sig_loopback =-5632;
8761: waveform_sig_loopback =-6183;
8762: waveform_sig_loopback =-6702;
8763: waveform_sig_loopback =-4526;
8764: waveform_sig_loopback =-6818;
8765: waveform_sig_loopback =-5892;
8766: waveform_sig_loopback =-5651;
8767: waveform_sig_loopback =-5682;
8768: waveform_sig_loopback =-6610;
8769: waveform_sig_loopback =-4952;
8770: waveform_sig_loopback =-5514;
8771: waveform_sig_loopback =-7084;
8772: waveform_sig_loopback =-4517;
8773: waveform_sig_loopback =-5810;
8774: waveform_sig_loopback =-6110;
8775: waveform_sig_loopback =-5619;
8776: waveform_sig_loopback =-4832;
8777: waveform_sig_loopback =-6024;
8778: waveform_sig_loopback =-6369;
8779: waveform_sig_loopback =-4135;
8780: waveform_sig_loopback =-5525;
8781: waveform_sig_loopback =-7012;
8782: waveform_sig_loopback =-4340;
8783: waveform_sig_loopback =-4421;
8784: waveform_sig_loopback =-6814;
8785: waveform_sig_loopback =-5560;
8786: waveform_sig_loopback =-3567;
8787: waveform_sig_loopback =-6513;
8788: waveform_sig_loopback =-4070;
8789: waveform_sig_loopback =-5304;
8790: waveform_sig_loopback =-8312;
8791: waveform_sig_loopback =-2269;
8792: waveform_sig_loopback =-4620;
8793: waveform_sig_loopback =-5891;
8794: waveform_sig_loopback =-5919;
8795: waveform_sig_loopback =-5298;
8796: waveform_sig_loopback =-2963;
8797: waveform_sig_loopback =-5291;
8798: waveform_sig_loopback =-6438;
8799: waveform_sig_loopback =-3573;
8800: waveform_sig_loopback =-5762;
8801: waveform_sig_loopback =-3929;
8802: waveform_sig_loopback =-5152;
8803: waveform_sig_loopback =-5443;
8804: waveform_sig_loopback =-3224;
8805: waveform_sig_loopback =-5837;
8806: waveform_sig_loopback =-4160;
8807: waveform_sig_loopback =-4432;
8808: waveform_sig_loopback =-4755;
8809: waveform_sig_loopback =-5013;
8810: waveform_sig_loopback =-3599;
8811: waveform_sig_loopback =-4439;
8812: waveform_sig_loopback =-5490;
8813: waveform_sig_loopback =-3414;
8814: waveform_sig_loopback =-4316;
8815: waveform_sig_loopback =-4705;
8816: waveform_sig_loopback =-4558;
8817: waveform_sig_loopback =-3135;
8818: waveform_sig_loopback =-4800;
8819: waveform_sig_loopback =-5031;
8820: waveform_sig_loopback =-2533;
8821: waveform_sig_loopback =-4410;
8822: waveform_sig_loopback =-5410;
8823: waveform_sig_loopback =-2804;
8824: waveform_sig_loopback =-3361;
8825: waveform_sig_loopback =-5153;
8826: waveform_sig_loopback =-4031;
8827: waveform_sig_loopback =-2324;
8828: waveform_sig_loopback =-4946;
8829: waveform_sig_loopback =-2572;
8830: waveform_sig_loopback =-4034;
8831: waveform_sig_loopback =-6557;
8832: waveform_sig_loopback =-896;
8833: waveform_sig_loopback =-3143;
8834: waveform_sig_loopback =-4311;
8835: waveform_sig_loopback =-4646;
8836: waveform_sig_loopback =-3430;
8837: waveform_sig_loopback =-1477;
8838: waveform_sig_loopback =-3981;
8839: waveform_sig_loopback =-4553;
8840: waveform_sig_loopback =-2279;
8841: waveform_sig_loopback =-3874;
8842: waveform_sig_loopback =-2342;
8843: waveform_sig_loopback =-4013;
8844: waveform_sig_loopback =-3393;
8845: waveform_sig_loopback =-1660;
8846: waveform_sig_loopback =-4466;
8847: waveform_sig_loopback =-2472;
8848: waveform_sig_loopback =-2984;
8849: waveform_sig_loopback =-2981;
8850: waveform_sig_loopback =-3243;
8851: waveform_sig_loopback =-2392;
8852: waveform_sig_loopback =-2593;
8853: waveform_sig_loopback =-3736;
8854: waveform_sig_loopback =-2012;
8855: waveform_sig_loopback =-2446;
8856: waveform_sig_loopback =-3367;
8857: waveform_sig_loopback =-2644;
8858: waveform_sig_loopback =-1396;
8859: waveform_sig_loopback =-3615;
8860: waveform_sig_loopback =-2907;
8861: waveform_sig_loopback =-890;
8862: waveform_sig_loopback =-3014;
8863: waveform_sig_loopback =-3509;
8864: waveform_sig_loopback =-1165;
8865: waveform_sig_loopback =-1647;
8866: waveform_sig_loopback =-3482;
8867: waveform_sig_loopback =-2374;
8868: waveform_sig_loopback =-494;
8869: waveform_sig_loopback =-3251;
8870: waveform_sig_loopback =-843;
8871: waveform_sig_loopback =-2478;
8872: waveform_sig_loopback =-4586;
8873: waveform_sig_loopback =797;
8874: waveform_sig_loopback =-1353;
8875: waveform_sig_loopback =-2656;
8876: waveform_sig_loopback =-2945;
8877: waveform_sig_loopback =-1283;
8878: waveform_sig_loopback =-92;
8879: waveform_sig_loopback =-2134;
8880: waveform_sig_loopback =-2549;
8881: waveform_sig_loopback =-845;
8882: waveform_sig_loopback =-1691;
8883: waveform_sig_loopback =-826;
8884: waveform_sig_loopback =-2278;
8885: waveform_sig_loopback =-1190;
8886: waveform_sig_loopback =-388;
8887: waveform_sig_loopback =-2283;
8888: waveform_sig_loopback =-701;
8889: waveform_sig_loopback =-1404;
8890: waveform_sig_loopback =-738;
8891: waveform_sig_loopback =-1824;
8892: waveform_sig_loopback =-307;
8893: waveform_sig_loopback =-741;
8894: waveform_sig_loopback =-2140;
8895: waveform_sig_loopback =177;
8896: waveform_sig_loopback =-797;
8897: waveform_sig_loopback =-1551;
8898: waveform_sig_loopback =-576;
8899: waveform_sig_loopback =289;
8900: waveform_sig_loopback =-1737;
8901: waveform_sig_loopback =-903;
8902: waveform_sig_loopback =906;
8903: waveform_sig_loopback =-1261;
8904: waveform_sig_loopback =-1421;
8905: waveform_sig_loopback =632;
8906: waveform_sig_loopback =165;
8907: waveform_sig_loopback =-1477;
8908: waveform_sig_loopback =-650;
8909: waveform_sig_loopback =1613;
8910: waveform_sig_loopback =-1530;
8911: waveform_sig_loopback =1044;
8912: waveform_sig_loopback =-514;
8913: waveform_sig_loopback =-2886;
8914: waveform_sig_loopback =2945;
8915: waveform_sig_loopback =471;
8916: waveform_sig_loopback =-1161;
8917: waveform_sig_loopback =-577;
8918: waveform_sig_loopback =414;
8919: waveform_sig_loopback =1679;
8920: waveform_sig_loopback =27;
8921: waveform_sig_loopback =-1060;
8922: waveform_sig_loopback =1376;
8923: waveform_sig_loopback =142;
8924: waveform_sig_loopback =781;
8925: waveform_sig_loopback =22;
8926: waveform_sig_loopback =429;
8927: waveform_sig_loopback =1486;
8928: waveform_sig_loopback =-221;
8929: waveform_sig_loopback =899;
8930: waveform_sig_loopback =774;
8931: waveform_sig_loopback =973;
8932: waveform_sig_loopback =29;
8933: waveform_sig_loopback =1845;
8934: waveform_sig_loopback =870;
8935: waveform_sig_loopback =-127;
8936: waveform_sig_loopback =2113;
8937: waveform_sig_loopback =1064;
8938: waveform_sig_loopback =316;
8939: waveform_sig_loopback =1499;
8940: waveform_sig_loopback =2075;
8941: waveform_sig_loopback =79;
8942: waveform_sig_loopback =1266;
8943: waveform_sig_loopback =2488;
8944: waveform_sig_loopback =752;
8945: waveform_sig_loopback =538;
8946: waveform_sig_loopback =2330;
8947: waveform_sig_loopback =2349;
8948: waveform_sig_loopback =9;
8949: waveform_sig_loopback =1458;
8950: waveform_sig_loopback =3658;
8951: waveform_sig_loopback =-217;
8952: waveform_sig_loopback =3536;
8953: waveform_sig_loopback =908;
8954: waveform_sig_loopback =-1004;
8955: waveform_sig_loopback =5349;
8956: waveform_sig_loopback =1668;
8957: waveform_sig_loopback =1013;
8958: waveform_sig_loopback =1377;
8959: waveform_sig_loopback =1987;
8960: waveform_sig_loopback =4037;
8961: waveform_sig_loopback =1389;
8962: waveform_sig_loopback =968;
8963: waveform_sig_loopback =3480;
8964: waveform_sig_loopback =1592;
8965: waveform_sig_loopback =2979;
8966: waveform_sig_loopback =1707;
8967: waveform_sig_loopback =2260;
8968: waveform_sig_loopback =3529;
8969: waveform_sig_loopback =1431;
8970: waveform_sig_loopback =2846;
8971: waveform_sig_loopback =2593;
8972: waveform_sig_loopback =2769;
8973: waveform_sig_loopback =1839;
8974: waveform_sig_loopback =3743;
8975: waveform_sig_loopback =2602;
8976: waveform_sig_loopback =1648;
8977: waveform_sig_loopback =4143;
8978: waveform_sig_loopback =2536;
8979: waveform_sig_loopback =2257;
8980: waveform_sig_loopback =3482;
8981: waveform_sig_loopback =3427;
8982: waveform_sig_loopback =2289;
8983: waveform_sig_loopback =2804;
8984: waveform_sig_loopback =4330;
8985: waveform_sig_loopback =2756;
8986: waveform_sig_loopback =1831;
8987: waveform_sig_loopback =4674;
8988: waveform_sig_loopback =3838;
8989: waveform_sig_loopback =1563;
8990: waveform_sig_loopback =3854;
8991: waveform_sig_loopback =4800;
8992: waveform_sig_loopback =1831;
8993: waveform_sig_loopback =5508;
8994: waveform_sig_loopback =1987;
8995: waveform_sig_loopback =1495;
8996: waveform_sig_loopback =6751;
8997: waveform_sig_loopback =3328;
8998: waveform_sig_loopback =3098;
8999: waveform_sig_loopback =2601;
9000: waveform_sig_loopback =4141;
9001: waveform_sig_loopback =5684;
9002: waveform_sig_loopback =2825;
9003: waveform_sig_loopback =2950;
9004: waveform_sig_loopback =4957;
9005: waveform_sig_loopback =3402;
9006: waveform_sig_loopback =4721;
9007: waveform_sig_loopback =3179;
9008: waveform_sig_loopback =4076;
9009: waveform_sig_loopback =5217;
9010: waveform_sig_loopback =3083;
9011: waveform_sig_loopback =4417;
9012: waveform_sig_loopback =4447;
9013: waveform_sig_loopback =4193;
9014: waveform_sig_loopback =3594;
9015: waveform_sig_loopback =5591;
9016: waveform_sig_loopback =3635;
9017: waveform_sig_loopback =3936;
9018: waveform_sig_loopback =5424;
9019: waveform_sig_loopback =4048;
9020: waveform_sig_loopback =4197;
9021: waveform_sig_loopback =4544;
9022: waveform_sig_loopback =5586;
9023: waveform_sig_loopback =3508;
9024: waveform_sig_loopback =4311;
9025: waveform_sig_loopback =6309;
9026: waveform_sig_loopback =3778;
9027: waveform_sig_loopback =3725;
9028: waveform_sig_loopback =6291;
9029: waveform_sig_loopback =5119;
9030: waveform_sig_loopback =3349;
9031: waveform_sig_loopback =5362;
9032: waveform_sig_loopback =6181;
9033: waveform_sig_loopback =3569;
9034: waveform_sig_loopback =6959;
9035: waveform_sig_loopback =3244;
9036: waveform_sig_loopback =3327;
9037: waveform_sig_loopback =8097;
9038: waveform_sig_loopback =4828;
9039: waveform_sig_loopback =4529;
9040: waveform_sig_loopback =3970;
9041: waveform_sig_loopback =5840;
9042: waveform_sig_loopback =7009;
9043: waveform_sig_loopback =4093;
9044: waveform_sig_loopback =4642;
9045: waveform_sig_loopback =6262;
9046: waveform_sig_loopback =4776;
9047: waveform_sig_loopback =6304;
9048: waveform_sig_loopback =4319;
9049: waveform_sig_loopback =5740;
9050: waveform_sig_loopback =6535;
9051: waveform_sig_loopback =4224;
9052: waveform_sig_loopback =6153;
9053: waveform_sig_loopback =5634;
9054: waveform_sig_loopback =5412;
9055: waveform_sig_loopback =5330;
9056: waveform_sig_loopback =6532;
9057: waveform_sig_loopback =5182;
9058: waveform_sig_loopback =5351;
9059: waveform_sig_loopback =6355;
9060: waveform_sig_loopback =5891;
9061: waveform_sig_loopback =5072;
9062: waveform_sig_loopback =6075;
9063: waveform_sig_loopback =6959;
9064: waveform_sig_loopback =4332;
9065: waveform_sig_loopback =6166;
9066: waveform_sig_loopback =7245;
9067: waveform_sig_loopback =4938;
9068: waveform_sig_loopback =5269;
9069: waveform_sig_loopback =7291;
9070: waveform_sig_loopback =6360;
9071: waveform_sig_loopback =4535;
9072: waveform_sig_loopback =6659;
9073: waveform_sig_loopback =7293;
9074: waveform_sig_loopback =4794;
9075: waveform_sig_loopback =8106;
9076: waveform_sig_loopback =4145;
9077: waveform_sig_loopback =4886;
9078: waveform_sig_loopback =8992;
9079: waveform_sig_loopback =6021;
9080: waveform_sig_loopback =5553;
9081: waveform_sig_loopback =5054;
9082: waveform_sig_loopback =7344;
9083: waveform_sig_loopback =7693;
9084: waveform_sig_loopback =5284;
9085: waveform_sig_loopback =5953;
9086: waveform_sig_loopback =6981;
9087: waveform_sig_loopback =6190;
9088: waveform_sig_loopback =7119;
9089: waveform_sig_loopback =5294;
9090: waveform_sig_loopback =7183;
9091: waveform_sig_loopback =7065;
9092: waveform_sig_loopback =5505;
9093: waveform_sig_loopback =7272;
9094: waveform_sig_loopback =6313;
9095: waveform_sig_loopback =6752;
9096: waveform_sig_loopback =6000;
9097: waveform_sig_loopback =7651;
9098: waveform_sig_loopback =6260;
9099: waveform_sig_loopback =6037;
9100: waveform_sig_loopback =7574;
9101: waveform_sig_loopback =6694;
9102: waveform_sig_loopback =5921;
9103: waveform_sig_loopback =7196;
9104: waveform_sig_loopback =7684;
9105: waveform_sig_loopback =5218;
9106: waveform_sig_loopback =7274;
9107: waveform_sig_loopback =7974;
9108: waveform_sig_loopback =5738;
9109: waveform_sig_loopback =6305;
9110: waveform_sig_loopback =8011;
9111: waveform_sig_loopback =7143;
9112: waveform_sig_loopback =5431;
9113: waveform_sig_loopback =7381;
9114: waveform_sig_loopback =8184;
9115: waveform_sig_loopback =5475;
9116: waveform_sig_loopback =8824;
9117: waveform_sig_loopback =5058;
9118: waveform_sig_loopback =5491;
9119: waveform_sig_loopback =9864;
9120: waveform_sig_loopback =6843;
9121: waveform_sig_loopback =5932;
9122: waveform_sig_loopback =6191;
9123: waveform_sig_loopback =7782;
9124: waveform_sig_loopback =8340;
9125: waveform_sig_loopback =6180;
9126: waveform_sig_loopback =6311;
9127: waveform_sig_loopback =7886;
9128: waveform_sig_loopback =6857;
9129: waveform_sig_loopback =7573;
9130: waveform_sig_loopback =6143;
9131: waveform_sig_loopback =7679;
9132: waveform_sig_loopback =7588;
9133: waveform_sig_loopback =6343;
9134: waveform_sig_loopback =7549;
9135: waveform_sig_loopback =6997;
9136: waveform_sig_loopback =7372;
9137: waveform_sig_loopback =6403;
9138: waveform_sig_loopback =8286;
9139: waveform_sig_loopback =6583;
9140: waveform_sig_loopback =6465;
9141: waveform_sig_loopback =8274;
9142: waveform_sig_loopback =6920;
9143: waveform_sig_loopback =6359;
9144: waveform_sig_loopback =7942;
9145: waveform_sig_loopback =7603;
9146: waveform_sig_loopback =5892;
9147: waveform_sig_loopback =7716;
9148: waveform_sig_loopback =8145;
9149: waveform_sig_loopback =6179;
9150: waveform_sig_loopback =6434;
9151: waveform_sig_loopback =8595;
9152: waveform_sig_loopback =7547;
9153: waveform_sig_loopback =5431;
9154: waveform_sig_loopback =7777;
9155: waveform_sig_loopback =8658;
9156: waveform_sig_loopback =5657;
9157: waveform_sig_loopback =9304;
9158: waveform_sig_loopback =4892;
9159: waveform_sig_loopback =6054;
9160: waveform_sig_loopback =10493;
9161: waveform_sig_loopback =6440;
9162: waveform_sig_loopback =6296;
9163: waveform_sig_loopback =6641;
9164: waveform_sig_loopback =7812;
9165: waveform_sig_loopback =8710;
9166: waveform_sig_loopback =6057;
9167: waveform_sig_loopback =6623;
9168: waveform_sig_loopback =8237;
9169: waveform_sig_loopback =6589;
9170: waveform_sig_loopback =7780;
9171: waveform_sig_loopback =6436;
9172: waveform_sig_loopback =7631;
9173: waveform_sig_loopback =7654;
9174: waveform_sig_loopback =6358;
9175: waveform_sig_loopback =7581;
9176: waveform_sig_loopback =7262;
9177: waveform_sig_loopback =7145;
9178: waveform_sig_loopback =6421;
9179: waveform_sig_loopback =8608;
9180: waveform_sig_loopback =6250;
9181: waveform_sig_loopback =6642;
9182: waveform_sig_loopback =8369;
9183: waveform_sig_loopback =6561;
9184: waveform_sig_loopback =6620;
9185: waveform_sig_loopback =7809;
9186: waveform_sig_loopback =7433;
9187: waveform_sig_loopback =6114;
9188: waveform_sig_loopback =7359;
9189: waveform_sig_loopback =8113;
9190: waveform_sig_loopback =6205;
9191: waveform_sig_loopback =6274;
9192: waveform_sig_loopback =8587;
9193: waveform_sig_loopback =7124;
9194: waveform_sig_loopback =5335;
9195: waveform_sig_loopback =8133;
9196: waveform_sig_loopback =7903;
9197: waveform_sig_loopback =5560;
9198: waveform_sig_loopback =9381;
9199: waveform_sig_loopback =4307;
9200: waveform_sig_loopback =6154;
9201: waveform_sig_loopback =10022;
9202: waveform_sig_loopback =6124;
9203: waveform_sig_loopback =6288;
9204: waveform_sig_loopback =6060;
9205: waveform_sig_loopback =7550;
9206: waveform_sig_loopback =8677;
9207: waveform_sig_loopback =5369;
9208: waveform_sig_loopback =6460;
9209: waveform_sig_loopback =7874;
9210: waveform_sig_loopback =6167;
9211: waveform_sig_loopback =7726;
9212: waveform_sig_loopback =5684;
9213: waveform_sig_loopback =7406;
9214: waveform_sig_loopback =7502;
9215: waveform_sig_loopback =5766;
9216: waveform_sig_loopback =7250;
9217: waveform_sig_loopback =6854;
9218: waveform_sig_loopback =6552;
9219: waveform_sig_loopback =6305;
9220: waveform_sig_loopback =8039;
9221: waveform_sig_loopback =5605;
9222: waveform_sig_loopback =6609;
9223: waveform_sig_loopback =7550;
9224: waveform_sig_loopback =6144;
9225: waveform_sig_loopback =6236;
9226: waveform_sig_loopback =7152;
9227: waveform_sig_loopback =7101;
9228: waveform_sig_loopback =5403;
9229: waveform_sig_loopback =6852;
9230: waveform_sig_loopback =7704;
9231: waveform_sig_loopback =5406;
9232: waveform_sig_loopback =5765;
9233: waveform_sig_loopback =8166;
9234: waveform_sig_loopback =6284;
9235: waveform_sig_loopback =4816;
9236: waveform_sig_loopback =7687;
9237: waveform_sig_loopback =6853;
9238: waveform_sig_loopback =5228;
9239: waveform_sig_loopback =8555;
9240: waveform_sig_loopback =3260;
9241: waveform_sig_loopback =6086;
9242: waveform_sig_loopback =8912;
9243: waveform_sig_loopback =5485;
9244: waveform_sig_loopback =5652;
9245: waveform_sig_loopback =5041;
9246: waveform_sig_loopback =7230;
9247: waveform_sig_loopback =7642;
9248: waveform_sig_loopback =4429;
9249: waveform_sig_loopback =6109;
9250: waveform_sig_loopback =6664;
9251: waveform_sig_loopback =5524;
9252: waveform_sig_loopback =6925;
9253: waveform_sig_loopback =4518;
9254: waveform_sig_loopback =6990;
9255: waveform_sig_loopback =6306;
9256: waveform_sig_loopback =4872;
9257: waveform_sig_loopback =6618;
9258: waveform_sig_loopback =5783;
9259: waveform_sig_loopback =5669;
9260: waveform_sig_loopback =5458;
9261: waveform_sig_loopback =6921;
9262: waveform_sig_loopback =4707;
9263: waveform_sig_loopback =5781;
9264: waveform_sig_loopback =6394;
9265: waveform_sig_loopback =5345;
9266: waveform_sig_loopback =5203;
9267: waveform_sig_loopback =6023;
9268: waveform_sig_loopback =6272;
9269: waveform_sig_loopback =4137;
9270: waveform_sig_loopback =6030;
9271: waveform_sig_loopback =6775;
9272: waveform_sig_loopback =3960;
9273: waveform_sig_loopback =5179;
9274: waveform_sig_loopback =6964;
9275: waveform_sig_loopback =4920;
9276: waveform_sig_loopback =4103;
9277: waveform_sig_loopback =6348;
9278: waveform_sig_loopback =5830;
9279: waveform_sig_loopback =4315;
9280: waveform_sig_loopback =7140;
9281: waveform_sig_loopback =2324;
9282: waveform_sig_loopback =5046;
9283: waveform_sig_loopback =7585;
9284: waveform_sig_loopback =4498;
9285: waveform_sig_loopback =4283;
9286: waveform_sig_loopback =4024;
9287: waveform_sig_loopback =6216;
9288: waveform_sig_loopback =6172;
9289: waveform_sig_loopback =3356;
9290: waveform_sig_loopback =5004;
9291: waveform_sig_loopback =5227;
9292: waveform_sig_loopback =4592;
9293: waveform_sig_loopback =5512;
9294: waveform_sig_loopback =3281;
9295: waveform_sig_loopback =5958;
9296: waveform_sig_loopback =4689;
9297: waveform_sig_loopback =3778;
9298: waveform_sig_loopback =5382;
9299: waveform_sig_loopback =4220;
9300: waveform_sig_loopback =4572;
9301: waveform_sig_loopback =4126;
9302: waveform_sig_loopback =5470;
9303: waveform_sig_loopback =3574;
9304: waveform_sig_loopback =4239;
9305: waveform_sig_loopback =5137;
9306: waveform_sig_loopback =4044;
9307: waveform_sig_loopback =3589;
9308: waveform_sig_loopback =4992;
9309: waveform_sig_loopback =4655;
9310: waveform_sig_loopback =2635;
9311: waveform_sig_loopback =4949;
9312: waveform_sig_loopback =5089;
9313: waveform_sig_loopback =2517;
9314: waveform_sig_loopback =4017;
9315: waveform_sig_loopback =5248;
9316: waveform_sig_loopback =3612;
9317: waveform_sig_loopback =2652;
9318: waveform_sig_loopback =4784;
9319: waveform_sig_loopback =4537;
9320: waveform_sig_loopback =2661;
9321: waveform_sig_loopback =5720;
9322: waveform_sig_loopback =796;
9323: waveform_sig_loopback =3569;
9324: waveform_sig_loopback =6222;
9325: waveform_sig_loopback =2826;
9326: waveform_sig_loopback =2626;
9327: waveform_sig_loopback =2769;
9328: waveform_sig_loopback =4632;
9329: waveform_sig_loopback =4471;
9330: waveform_sig_loopback =1953;
9331: waveform_sig_loopback =3404;
9332: waveform_sig_loopback =3666;
9333: waveform_sig_loopback =3160;
9334: waveform_sig_loopback =3639;
9335: waveform_sig_loopback =1965;
9336: waveform_sig_loopback =4391;
9337: waveform_sig_loopback =2821;
9338: waveform_sig_loopback =2545;
9339: waveform_sig_loopback =3499;
9340: waveform_sig_loopback =2688;
9341: waveform_sig_loopback =3131;
9342: waveform_sig_loopback =2190;
9343: waveform_sig_loopback =4178;
9344: waveform_sig_loopback =1782;
9345: waveform_sig_loopback =2460;
9346: waveform_sig_loopback =3834;
9347: waveform_sig_loopback =1992;
9348: waveform_sig_loopback =2200;
9349: waveform_sig_loopback =3353;
9350: waveform_sig_loopback =2708;
9351: waveform_sig_loopback =1254;
9352: waveform_sig_loopback =3236;
9353: waveform_sig_loopback =3282;
9354: waveform_sig_loopback =868;
9355: waveform_sig_loopback =2385;
9356: waveform_sig_loopback =3470;
9357: waveform_sig_loopback =1958;
9358: waveform_sig_loopback =871;
9359: waveform_sig_loopback =3182;
9360: waveform_sig_loopback =2808;
9361: waveform_sig_loopback =820;
9362: waveform_sig_loopback =4118;
9363: waveform_sig_loopback =-1130;
9364: waveform_sig_loopback =1910;
9365: waveform_sig_loopback =4582;
9366: waveform_sig_loopback =863;
9367: waveform_sig_loopback =817;
9368: waveform_sig_loopback =1246;
9369: waveform_sig_loopback =2621;
9370: waveform_sig_loopback =2835;
9371: waveform_sig_loopback =150;
9372: waveform_sig_loopback =1374;
9373: waveform_sig_loopback =2212;
9374: waveform_sig_loopback =1139;
9375: waveform_sig_loopback =1776;
9376: waveform_sig_loopback =446;
9377: waveform_sig_loopback =2202;
9378: waveform_sig_loopback =1305;
9379: waveform_sig_loopback =680;
9380: waveform_sig_loopback =1487;
9381: waveform_sig_loopback =1306;
9382: waveform_sig_loopback =911;
9383: waveform_sig_loopback =656;
9384: waveform_sig_loopback =2316;
9385: waveform_sig_loopback =-271;
9386: waveform_sig_loopback =992;
9387: waveform_sig_loopback =1758;
9388: waveform_sig_loopback =194;
9389: waveform_sig_loopback =327;
9390: waveform_sig_loopback =1702;
9391: waveform_sig_loopback =645;
9392: waveform_sig_loopback =-465;
9393: waveform_sig_loopback =1493;
9394: waveform_sig_loopback =1123;
9395: waveform_sig_loopback =-668;
9396: waveform_sig_loopback =291;
9397: waveform_sig_loopback =1788;
9398: waveform_sig_loopback =70;
9399: waveform_sig_loopback =-1313;
9400: waveform_sig_loopback =1876;
9401: waveform_sig_loopback =445;
9402: waveform_sig_loopback =-883;
9403: waveform_sig_loopback =2406;
9404: waveform_sig_loopback =-3543;
9405: waveform_sig_loopback =688;
9406: waveform_sig_loopback =2520;
9407: waveform_sig_loopback =-1357;
9408: waveform_sig_loopback =-595;
9409: waveform_sig_loopback =-909;
9410: waveform_sig_loopback =881;
9411: waveform_sig_loopback =1070;
9412: waveform_sig_loopback =-2168;
9413: waveform_sig_loopback =-10;
9414: waveform_sig_loopback =156;
9415: waveform_sig_loopback =-856;
9416: waveform_sig_loopback =192;
9417: waveform_sig_loopback =-1726;
9418: waveform_sig_loopback =539;
9419: waveform_sig_loopback =-647;
9420: waveform_sig_loopback =-1335;
9421: waveform_sig_loopback =-257;
9422: waveform_sig_loopback =-685;
9423: waveform_sig_loopback =-1154;
9424: waveform_sig_loopback =-1039;
9425: waveform_sig_loopback =358;
9426: waveform_sig_loopback =-2363;
9427: waveform_sig_loopback =-651;
9428: waveform_sig_loopback =-217;
9429: waveform_sig_loopback =-1801;
9430: waveform_sig_loopback =-1341;
9431: waveform_sig_loopback =-390;
9432: waveform_sig_loopback =-1260;
9433: waveform_sig_loopback =-2191;
9434: waveform_sig_loopback =-661;
9435: waveform_sig_loopback =-537;
9436: waveform_sig_loopback =-2655;
9437: waveform_sig_loopback =-1746;
9438: waveform_sig_loopback =269;
9439: waveform_sig_loopback =-2329;
9440: waveform_sig_loopback =-2890;
9441: waveform_sig_loopback =264;
9442: waveform_sig_loopback =-2035;
9443: waveform_sig_loopback =-2053;
9444: waveform_sig_loopback =89;
9445: waveform_sig_loopback =-5501;
9446: waveform_sig_loopback =-472;
9447: waveform_sig_loopback =-84;
9448: waveform_sig_loopback =-2739;
9449: waveform_sig_loopback =-2654;
9450: waveform_sig_loopback =-2946;
9451: waveform_sig_loopback =-452;
9452: waveform_sig_loopback =-1249;
9453: waveform_sig_loopback =-3904;
9454: waveform_sig_loopback =-1714;
9455: waveform_sig_loopback =-2000;
9456: waveform_sig_loopback =-2387;
9457: waveform_sig_loopback =-1876;
9458: waveform_sig_loopback =-3599;
9459: waveform_sig_loopback =-1131;
9460: waveform_sig_loopback =-2601;
9461: waveform_sig_loopback =-3133;
9462: waveform_sig_loopback =-2098;
9463: waveform_sig_loopback =-2414;
9464: waveform_sig_loopback =-3142;
9465: waveform_sig_loopback =-2597;
9466: waveform_sig_loopback =-1677;
9467: waveform_sig_loopback =-4235;
9468: waveform_sig_loopback =-2028;
9469: waveform_sig_loopback =-2617;
9470: waveform_sig_loopback =-3234;
9471: waveform_sig_loopback =-3209;
9472: waveform_sig_loopback =-2398;
9473: waveform_sig_loopback =-2609;
9474: waveform_sig_loopback =-4554;
9475: waveform_sig_loopback =-2020;
9476: waveform_sig_loopback =-2342;
9477: waveform_sig_loopback =-4904;
9478: waveform_sig_loopback =-2876;
9479: waveform_sig_loopback =-1902;
9480: waveform_sig_loopback =-4091;
9481: waveform_sig_loopback =-4396;
9482: waveform_sig_loopback =-1892;
9483: waveform_sig_loopback =-3623;
9484: waveform_sig_loopback =-3762;
9485: waveform_sig_loopback =-1956;
9486: waveform_sig_loopback =-7088;
9487: waveform_sig_loopback =-2248;
9488: waveform_sig_loopback =-1834;
9489: waveform_sig_loopback =-4466;
9490: waveform_sig_loopback =-4504;
9491: waveform_sig_loopback =-4552;
9492: waveform_sig_loopback =-2103;
9493: waveform_sig_loopback =-3142;
9494: waveform_sig_loopback =-5651;
9495: waveform_sig_loopback =-3207;
9496: waveform_sig_loopback =-3984;
9497: waveform_sig_loopback =-3921;
9498: waveform_sig_loopback =-3806;
9499: waveform_sig_loopback =-5288;
9500: waveform_sig_loopback =-2457;
9501: waveform_sig_loopback =-4668;
9502: waveform_sig_loopback =-4924;
9503: waveform_sig_loopback =-3469;
9504: waveform_sig_loopback =-4302;
9505: waveform_sig_loopback =-4653;
9506: waveform_sig_loopback =-4328;
9507: waveform_sig_loopback =-3683;
9508: waveform_sig_loopback =-5222;
9509: waveform_sig_loopback =-4184;
9510: waveform_sig_loopback =-4167;
9511: waveform_sig_loopback =-4643;
9512: waveform_sig_loopback =-5218;
9513: waveform_sig_loopback =-3492;
9514: waveform_sig_loopback =-4743;
9515: waveform_sig_loopback =-6008;
9516: waveform_sig_loopback =-3269;
9517: waveform_sig_loopback =-4443;
9518: waveform_sig_loopback =-6286;
9519: waveform_sig_loopback =-4348;
9520: waveform_sig_loopback =-3594;
9521: waveform_sig_loopback =-5640;
9522: waveform_sig_loopback =-6007;
9523: waveform_sig_loopback =-3314;
9524: waveform_sig_loopback =-5200;
9525: waveform_sig_loopback =-5249;
9526: waveform_sig_loopback =-3639;
9527: waveform_sig_loopback =-8501;
9528: waveform_sig_loopback =-3594;
9529: waveform_sig_loopback =-3510;
9530: waveform_sig_loopback =-5934;
9531: waveform_sig_loopback =-6164;
9532: waveform_sig_loopback =-5757;
9533: waveform_sig_loopback =-3593;
9534: waveform_sig_loopback =-4947;
9535: waveform_sig_loopback =-6782;
9536: waveform_sig_loopback =-4781;
9537: waveform_sig_loopback =-5512;
9538: waveform_sig_loopback =-5078;
9539: waveform_sig_loopback =-5435;
9540: waveform_sig_loopback =-6497;
9541: waveform_sig_loopback =-3956;
9542: waveform_sig_loopback =-6304;
9543: waveform_sig_loopback =-5675;
9544: waveform_sig_loopback =-5232;
9545: waveform_sig_loopback =-5757;
9546: waveform_sig_loopback =-5723;
9547: waveform_sig_loopback =-5908;
9548: waveform_sig_loopback =-4731;
9549: waveform_sig_loopback =-6906;
9550: waveform_sig_loopback =-5546;
9551: waveform_sig_loopback =-5082;
9552: waveform_sig_loopback =-6414;
9553: waveform_sig_loopback =-6361;
9554: waveform_sig_loopback =-4662;
9555: waveform_sig_loopback =-6311;
9556: waveform_sig_loopback =-7013;
9557: waveform_sig_loopback =-4695;
9558: waveform_sig_loopback =-5784;
9559: waveform_sig_loopback =-7331;
9560: waveform_sig_loopback =-5701;
9561: waveform_sig_loopback =-4866;
9562: waveform_sig_loopback =-6864;
9563: waveform_sig_loopback =-7188;
9564: waveform_sig_loopback =-4509;
9565: waveform_sig_loopback =-6488;
9566: waveform_sig_loopback =-6362;
9567: waveform_sig_loopback =-4912;
9568: waveform_sig_loopback =-9594;
9569: waveform_sig_loopback =-4847;
9570: waveform_sig_loopback =-4527;
9571: waveform_sig_loopback =-7158;
9572: waveform_sig_loopback =-7468;
9573: waveform_sig_loopback =-6487;
9574: waveform_sig_loopback =-5033;
9575: waveform_sig_loopback =-5862;
9576: waveform_sig_loopback =-7836;
9577: waveform_sig_loopback =-6112;
9578: waveform_sig_loopback =-6125;
9579: waveform_sig_loopback =-6421;
9580: waveform_sig_loopback =-6486;
9581: waveform_sig_loopback =-7277;
9582: waveform_sig_loopback =-5325;
9583: waveform_sig_loopback =-7104;
9584: waveform_sig_loopback =-6713;
9585: waveform_sig_loopback =-6432;
9586: waveform_sig_loopback =-6475;
9587: waveform_sig_loopback =-6949;
9588: waveform_sig_loopback =-6690;
9589: waveform_sig_loopback =-5647;
9590: waveform_sig_loopback =-8023;
9591: waveform_sig_loopback =-6220;
9592: waveform_sig_loopback =-6041;
9593: waveform_sig_loopback =-7471;
9594: waveform_sig_loopback =-7090;
9595: waveform_sig_loopback =-5572;
9596: waveform_sig_loopback =-7400;
9597: waveform_sig_loopback =-7613;
9598: waveform_sig_loopback =-5625;
9599: waveform_sig_loopback =-6764;
9600: waveform_sig_loopback =-7947;
9601: waveform_sig_loopback =-6707;
9602: waveform_sig_loopback =-5517;
9603: waveform_sig_loopback =-7691;
9604: waveform_sig_loopback =-8130;
9605: waveform_sig_loopback =-4908;
9606: waveform_sig_loopback =-7605;
9607: waveform_sig_loopback =-6923;
9608: waveform_sig_loopback =-5653;
9609: waveform_sig_loopback =-10624;
9610: waveform_sig_loopback =-5093;
9611: waveform_sig_loopback =-5416;
9612: waveform_sig_loopback =-8094;
9613: waveform_sig_loopback =-7892;
9614: waveform_sig_loopback =-7276;
9615: waveform_sig_loopback =-5739;
9616: waveform_sig_loopback =-6422;
9617: waveform_sig_loopback =-8760;
9618: waveform_sig_loopback =-6548;
9619: waveform_sig_loopback =-6789;
9620: waveform_sig_loopback =-7273;
9621: waveform_sig_loopback =-6913;
9622: waveform_sig_loopback =-7964;
9623: waveform_sig_loopback =-5976;
9624: waveform_sig_loopback =-7544;
9625: waveform_sig_loopback =-7463;
9626: waveform_sig_loopback =-6876;
9627: waveform_sig_loopback =-6949;
9628: waveform_sig_loopback =-7788;
9629: waveform_sig_loopback =-6897;
9630: waveform_sig_loopback =-6295;
9631: waveform_sig_loopback =-8668;
9632: waveform_sig_loopback =-6384;
9633: waveform_sig_loopback =-6768;
9634: waveform_sig_loopback =-7892;
9635: waveform_sig_loopback =-7298;
9636: waveform_sig_loopback =-6295;
9637: waveform_sig_loopback =-7641;
9638: waveform_sig_loopback =-7981;
9639: waveform_sig_loopback =-6135;
9640: waveform_sig_loopback =-6988;
9641: waveform_sig_loopback =-8519;
9642: waveform_sig_loopback =-6903;
9643: waveform_sig_loopback =-5811;
9644: waveform_sig_loopback =-8339;
9645: waveform_sig_loopback =-8221;
9646: waveform_sig_loopback =-5132;
9647: waveform_sig_loopback =-8240;
9648: waveform_sig_loopback =-6859;
9649: waveform_sig_loopback =-6167;
9650: waveform_sig_loopback =-11033;
9651: waveform_sig_loopback =-4892;
9652: waveform_sig_loopback =-6086;
9653: waveform_sig_loopback =-8279;
9654: waveform_sig_loopback =-7859;
9655: waveform_sig_loopback =-7838;
9656: waveform_sig_loopback =-5548;
9657: waveform_sig_loopback =-6823;
9658: waveform_sig_loopback =-9133;
9659: waveform_sig_loopback =-6207;
9660: waveform_sig_loopback =-7414;
9661: waveform_sig_loopback =-7109;
9662: waveform_sig_loopback =-7000;
9663: waveform_sig_loopback =-8303;
9664: waveform_sig_loopback =-5725;
9665: waveform_sig_loopback =-7892;
9666: waveform_sig_loopback =-7473;
9667: waveform_sig_loopback =-6812;
9668: waveform_sig_loopback =-7159;
9669: waveform_sig_loopback =-7784;
9670: waveform_sig_loopback =-6747;
9671: waveform_sig_loopback =-6548;
9672: waveform_sig_loopback =-8604;
9673: waveform_sig_loopback =-6245;
9674: waveform_sig_loopback =-6960;
9675: waveform_sig_loopback =-7734;
9676: waveform_sig_loopback =-7290;
9677: waveform_sig_loopback =-6381;
9678: waveform_sig_loopback =-7353;
9679: waveform_sig_loopback =-8089;
9680: waveform_sig_loopback =-6069;
9681: waveform_sig_loopback =-6772;
9682: waveform_sig_loopback =-8582;
9683: waveform_sig_loopback =-6472;
9684: waveform_sig_loopback =-5847;
9685: waveform_sig_loopback =-8397;
9686: waveform_sig_loopback =-7639;
9687: waveform_sig_loopback =-5189;
9688: waveform_sig_loopback =-8240;
9689: waveform_sig_loopback =-6298;
9690: waveform_sig_loopback =-6380;
9691: waveform_sig_loopback =-10635;
9692: waveform_sig_loopback =-4425;
9693: waveform_sig_loopback =-6220;
9694: waveform_sig_loopback =-7736;
9695: waveform_sig_loopback =-7751;
9696: waveform_sig_loopback =-7588;
9697: waveform_sig_loopback =-4828;
9698: waveform_sig_loopback =-6954;
9699: waveform_sig_loopback =-8602;
9700: waveform_sig_loopback =-5710;
9701: waveform_sig_loopback =-7448;
9702: waveform_sig_loopback =-6300;
9703: waveform_sig_loopback =-7017;
9704: waveform_sig_loopback =-7834;
9705: waveform_sig_loopback =-5133;
9706: waveform_sig_loopback =-7846;
9707: waveform_sig_loopback =-6802;
9708: waveform_sig_loopback =-6443;
9709: waveform_sig_loopback =-6823;
9710: waveform_sig_loopback =-7215;
9711: waveform_sig_loopback =-6294;
9712: waveform_sig_loopback =-6272;
9713: waveform_sig_loopback =-7937;
9714: waveform_sig_loopback =-5751;
9715: waveform_sig_loopback =-6698;
9716: waveform_sig_loopback =-7007;
9717: waveform_sig_loopback =-6777;
9718: waveform_sig_loopback =-5875;
9719: waveform_sig_loopback =-6756;
9720: waveform_sig_loopback =-7722;
9721: waveform_sig_loopback =-5047;
9722: waveform_sig_loopback =-6425;
9723: waveform_sig_loopback =-8326;
9724: waveform_sig_loopback =-5220;
9725: waveform_sig_loopback =-5782;
9726: waveform_sig_loopback =-7596;
9727: waveform_sig_loopback =-6767;
9728: waveform_sig_loopback =-4962;
9729: waveform_sig_loopback =-7131;
9730: waveform_sig_loopback =-5703;
9731: waveform_sig_loopback =-6003;
9732: waveform_sig_loopback =-9423;
9733: waveform_sig_loopback =-4001;
9734: waveform_sig_loopback =-5367;
9735: waveform_sig_loopback =-6959;
9736: waveform_sig_loopback =-7370;
9737: waveform_sig_loopback =-6321;
9738: waveform_sig_loopback =-4311;
9739: waveform_sig_loopback =-6349;
9740: waveform_sig_loopback =-7460;
9741: waveform_sig_loopback =-5207;
9742: waveform_sig_loopback =-6558;
9743: waveform_sig_loopback =-5339;
9744: waveform_sig_loopback =-6445;
9745: waveform_sig_loopback =-6746;
9746: waveform_sig_loopback =-4340;
9747: waveform_sig_loopback =-7137;
9748: waveform_sig_loopback =-5663;
9749: waveform_sig_loopback =-5715;
9750: waveform_sig_loopback =-6049;
9751: waveform_sig_loopback =-6020;
9752: waveform_sig_loopback =-5524;
9753: waveform_sig_loopback =-5447;
9754: waveform_sig_loopback =-6696;
9755: waveform_sig_loopback =-5180;
9756: waveform_sig_loopback =-5373;
9757: waveform_sig_loopback =-6165;
9758: waveform_sig_loopback =-6057;
9759: waveform_sig_loopback =-4286;
9760: waveform_sig_loopback =-6398;
9761: waveform_sig_loopback =-6414;
9762: waveform_sig_loopback =-3828;
9763: waveform_sig_loopback =-5950;
9764: waveform_sig_loopback =-6687;
9765: waveform_sig_loopback =-4437;
9766: waveform_sig_loopback =-4752;
9767: waveform_sig_loopback =-6276;
9768: waveform_sig_loopback =-5963;
9769: waveform_sig_loopback =-3633;
9770: waveform_sig_loopback =-6102;
9771: waveform_sig_loopback =-4664;
9772: waveform_sig_loopback =-4846;
9773: waveform_sig_loopback =-8326;
9774: waveform_sig_loopback =-2756;
9775: waveform_sig_loopback =-4150;
9776: waveform_sig_loopback =-6028;
9777: waveform_sig_loopback =-6118;
9778: waveform_sig_loopback =-4887;
9779: waveform_sig_loopback =-3392;
9780: waveform_sig_loopback =-5141;
9781: waveform_sig_loopback =-6127;
9782: waveform_sig_loopback =-4138;
9783: waveform_sig_loopback =-5143;
9784: waveform_sig_loopback =-4193;
9785: waveform_sig_loopback =-5371;
9786: waveform_sig_loopback =-5032;
9787: waveform_sig_loopback =-3492;
9788: waveform_sig_loopback =-5778;
9789: waveform_sig_loopback =-4107;
9790: waveform_sig_loopback =-4699;
9791: waveform_sig_loopback =-4441;
9792: waveform_sig_loopback =-4854;
9793: waveform_sig_loopback =-4300;
9794: waveform_sig_loopback =-3721;
9795: waveform_sig_loopback =-5668;
9796: waveform_sig_loopback =-3685;
9797: waveform_sig_loopback =-3812;
9798: waveform_sig_loopback =-5228;
9799: waveform_sig_loopback =-4116;
9800: waveform_sig_loopback =-3116;
9801: waveform_sig_loopback =-5196;
9802: waveform_sig_loopback =-4516;
9803: waveform_sig_loopback =-2770;
9804: waveform_sig_loopback =-4457;
9805: waveform_sig_loopback =-5095;
9806: waveform_sig_loopback =-3198;
9807: waveform_sig_loopback =-3110;
9808: waveform_sig_loopback =-4964;
9809: waveform_sig_loopback =-4528;
9810: waveform_sig_loopback =-1892;
9811: waveform_sig_loopback =-4902;
9812: waveform_sig_loopback =-2983;
9813: waveform_sig_loopback =-3411;
9814: waveform_sig_loopback =-6930;
9815: waveform_sig_loopback =-1003;
9816: waveform_sig_loopback =-2711;
9817: waveform_sig_loopback =-4716;
9818: waveform_sig_loopback =-4365;
9819: waveform_sig_loopback =-3284;
9820: waveform_sig_loopback =-2014;
9821: waveform_sig_loopback =-3356;
9822: waveform_sig_loopback =-4745;
9823: waveform_sig_loopback =-2554;
9824: waveform_sig_loopback =-3262;
9825: waveform_sig_loopback =-3010;
9826: waveform_sig_loopback =-3550;
9827: waveform_sig_loopback =-3347;
9828: waveform_sig_loopback =-2231;
9829: waveform_sig_loopback =-3705;
9830: waveform_sig_loopback =-2887;
9831: waveform_sig_loopback =-3077;
9832: waveform_sig_loopback =-2453;
9833: waveform_sig_loopback =-3755;
9834: waveform_sig_loopback =-2121;
9835: waveform_sig_loopback =-2390;
9836: waveform_sig_loopback =-4141;
9837: waveform_sig_loopback =-1548;
9838: waveform_sig_loopback =-2594;
9839: waveform_sig_loopback =-3392;
9840: waveform_sig_loopback =-2323;
9841: waveform_sig_loopback =-1738;
9842: waveform_sig_loopback =-3387;
9843: waveform_sig_loopback =-2795;
9844: waveform_sig_loopback =-1174;
9845: waveform_sig_loopback =-2831;
9846: waveform_sig_loopback =-3488;
9847: waveform_sig_loopback =-1387;
9848: waveform_sig_loopback =-1233;
9849: waveform_sig_loopback =-3545;
9850: waveform_sig_loopback =-2909;
9851: waveform_sig_loopback =287;
9852: waveform_sig_loopback =-3562;
9853: waveform_sig_loopback =-1000;
9854: waveform_sig_loopback =-1933;
9855: waveform_sig_loopback =-5343;
9856: waveform_sig_loopback =1471;
9857: waveform_sig_loopback =-1597;
9858: waveform_sig_loopback =-3012;
9859: waveform_sig_loopback =-2148;
9860: waveform_sig_loopback =-2021;
9861: waveform_sig_loopback =94;
9862: waveform_sig_loopback =-1835;
9863: waveform_sig_loopback =-3136;
9864: waveform_sig_loopback =-246;
9865: waveform_sig_loopback =-2086;
9866: waveform_sig_loopback =-1092;
9867: waveform_sig_loopback =-1600;
9868: waveform_sig_loopback =-1888;
9869: waveform_sig_loopback =-190;
9870: waveform_sig_loopback =-2087;
9871: waveform_sig_loopback =-1082;
9872: waveform_sig_loopback =-1037;
9873: waveform_sig_loopback =-940;
9874: waveform_sig_loopback =-1908;
9875: waveform_sig_loopback =-76;
9876: waveform_sig_loopback =-833;
9877: waveform_sig_loopback =-2269;
9878: waveform_sig_loopback =421;
9879: waveform_sig_loopback =-1002;
9880: waveform_sig_loopback =-1456;
9881: waveform_sig_loopback =-376;
9882: waveform_sig_loopback =-134;
9883: waveform_sig_loopback =-1261;
9884: waveform_sig_loopback =-1061;
9885: waveform_sig_loopback =571;
9886: waveform_sig_loopback =-594;
9887: waveform_sig_loopback =-1914;
9888: waveform_sig_loopback =641;
9889: waveform_sig_loopback =600;
9890: waveform_sig_loopback =-2017;
9891: waveform_sig_loopback =-278;
9892: waveform_sig_loopback =1510;
9893: waveform_sig_loopback =-1864;
9894: waveform_sig_loopback =1562;
9895: waveform_sig_loopback =-814;
9896: waveform_sig_loopback =-3007;
9897: waveform_sig_loopback =3226;
9898: waveform_sig_loopback =-42;
9899: waveform_sig_loopback =-579;
9900: waveform_sig_loopback =-829;
9901: waveform_sig_loopback =29;
9902: waveform_sig_loopback =2336;
9903: waveform_sig_loopback =-458;
9904: waveform_sig_loopback =-946;
9905: waveform_sig_loopback =1586;
9906: waveform_sig_loopback =-263;
9907: waveform_sig_loopback =1176;
9908: waveform_sig_loopback =-95;
9909: waveform_sig_loopback =189;
9910: waveform_sig_loopback =1938;
9911: waveform_sig_loopback =-376;
9912: waveform_sig_loopback =848;
9913: waveform_sig_loopback =946;
9914: waveform_sig_loopback =866;
9915: waveform_sig_loopback =40;
9916: waveform_sig_loopback =1971;
9917: waveform_sig_loopback =591;
9918: waveform_sig_loopback =115;
9919: waveform_sig_loopback =2168;
9920: waveform_sig_loopback =596;
9921: waveform_sig_loopback =909;
9922: waveform_sig_loopback =1059;
9923: waveform_sig_loopback =2049;
9924: waveform_sig_loopback =583;
9925: waveform_sig_loopback =538;
9926: waveform_sig_loopback =2993;
9927: waveform_sig_loopback =833;
9928: waveform_sig_loopback =15;
9929: waveform_sig_loopback =2898;
9930: waveform_sig_loopback =2002;
9931: waveform_sig_loopback =79;
9932: waveform_sig_loopback =1742;
9933: waveform_sig_loopback =3038;
9934: waveform_sig_loopback =395;
9935: waveform_sig_loopback =3339;
9936: waveform_sig_loopback =716;
9937: waveform_sig_loopback =-547;
9938: waveform_sig_loopback =4781;
9939: waveform_sig_loopback =1949;
9940: waveform_sig_loopback =1334;
9941: waveform_sig_loopback =808;
9942: waveform_sig_loopback =2342;
9943: waveform_sig_loopback =3959;
9944: waveform_sig_loopback =1325;
9945: waveform_sig_loopback =1157;
9946: waveform_sig_loopback =3320;
9947: waveform_sig_loopback =1581;
9948: waveform_sig_loopback =3211;
9949: waveform_sig_loopback =1511;
9950: waveform_sig_loopback =2166;
9951: waveform_sig_loopback =3872;
9952: waveform_sig_loopback =1115;
9953: waveform_sig_loopback =2998;
9954: waveform_sig_loopback =2729;
9955: waveform_sig_loopback =2351;
9956: waveform_sig_loopback =2383;
9957: waveform_sig_loopback =3408;
9958: waveform_sig_loopback =2439;
9959: waveform_sig_loopback =2257;
9960: waveform_sig_loopback =3365;
9961: waveform_sig_loopback =3011;
9962: waveform_sig_loopback =2325;
9963: waveform_sig_loopback =2802;
9964: waveform_sig_loopback =4298;
9965: waveform_sig_loopback =1657;
9966: waveform_sig_loopback =2900;
9967: waveform_sig_loopback =4642;
9968: waveform_sig_loopback =2280;
9969: waveform_sig_loopback =2252;
9970: waveform_sig_loopback =4389;
9971: waveform_sig_loopback =3848;
9972: waveform_sig_loopback =1869;
9973: waveform_sig_loopback =3522;
9974: waveform_sig_loopback =4822;
9975: waveform_sig_loopback =2123;
9976: waveform_sig_loopback =5176;
9977: waveform_sig_loopback =2250;
9978: waveform_sig_loopback =1516;
9979: waveform_sig_loopback =6376;
9980: waveform_sig_loopback =3722;
9981: waveform_sig_loopback =3008;
9982: waveform_sig_loopback =2372;
9983: waveform_sig_loopback =4514;
9984: waveform_sig_loopback =5300;
9985: waveform_sig_loopback =2981;
9986: waveform_sig_loopback =3199;
9987: waveform_sig_loopback =4612;
9988: waveform_sig_loopback =3613;
9989: waveform_sig_loopback =4723;
9990: waveform_sig_loopback =2978;
9991: waveform_sig_loopback =4360;
9992: waveform_sig_loopback =5042;
9993: waveform_sig_loopback =2900;
9994: waveform_sig_loopback =4895;
9995: waveform_sig_loopback =3968;
9996: waveform_sig_loopback =4397;
9997: waveform_sig_loopback =3782;
9998: waveform_sig_loopback =4929;
9999: waveform_sig_loopback =4408;
10000: waveform_sig_loopback =3490;
10001: waveform_sig_loopback =5204;
10002: waveform_sig_loopback =4677;
10003: waveform_sig_loopback =3602;
10004: waveform_sig_loopback =4867;
10005: waveform_sig_loopback =5592;
10006: waveform_sig_loopback =3205;
10007: waveform_sig_loopback =4753;
10008: waveform_sig_loopback =5951;
10009: waveform_sig_loopback =3847;
10010: waveform_sig_loopback =3992;
10011: waveform_sig_loopback =5934;
10012: waveform_sig_loopback =5332;
10013: waveform_sig_loopback =3518;
10014: waveform_sig_loopback =5019;
10015: waveform_sig_loopback =6487;
10016: waveform_sig_loopback =3597;
10017: waveform_sig_loopback =6582;
10018: waveform_sig_loopback =3858;
10019: waveform_sig_loopback =2949;
10020: waveform_sig_loopback =7906;
10021: waveform_sig_loopback =5335;
10022: waveform_sig_loopback =4081;
10023: waveform_sig_loopback =4185;
10024: waveform_sig_loopback =5972;
10025: waveform_sig_loopback =6485;
10026: waveform_sig_loopback =4767;
10027: waveform_sig_loopback =4346;
10028: waveform_sig_loopback =6043;
10029: waveform_sig_loopback =5259;
10030: waveform_sig_loopback =5767;
10031: waveform_sig_loopback =4648;
10032: waveform_sig_loopback =5764;
10033: waveform_sig_loopback =6112;
10034: waveform_sig_loopback =4750;
10035: waveform_sig_loopback =5889;
10036: waveform_sig_loopback =5388;
10037: waveform_sig_loopback =5980;
10038: waveform_sig_loopback =4781;
10039: waveform_sig_loopback =6700;
10040: waveform_sig_loopback =5472;
10041: waveform_sig_loopback =4751;
10042: waveform_sig_loopback =6866;
10043: waveform_sig_loopback =5659;
10044: waveform_sig_loopback =4997;
10045: waveform_sig_loopback =6340;
10046: waveform_sig_loopback =6614;
10047: waveform_sig_loopback =4575;
10048: waveform_sig_loopback =6166;
10049: waveform_sig_loopback =7000;
10050: waveform_sig_loopback =5192;
10051: waveform_sig_loopback =5268;
10052: waveform_sig_loopback =6975;
10053: waveform_sig_loopback =6680;
10054: waveform_sig_loopback =4516;
10055: waveform_sig_loopback =6263;
10056: waveform_sig_loopback =7849;
10057: waveform_sig_loopback =4378;
10058: waveform_sig_loopback =8074;
10059: waveform_sig_loopback =4836;
10060: waveform_sig_loopback =3955;
10061: waveform_sig_loopback =9555;
10062: waveform_sig_loopback =6026;
10063: waveform_sig_loopback =5205;
10064: waveform_sig_loopback =5733;
10065: waveform_sig_loopback =6603;
10066: waveform_sig_loopback =7974;
10067: waveform_sig_loopback =5675;
10068: waveform_sig_loopback =5265;
10069: waveform_sig_loopback =7577;
10070: waveform_sig_loopback =5911;
10071: waveform_sig_loopback =6970;
10072: waveform_sig_loopback =5863;
10073: waveform_sig_loopback =6550;
10074: waveform_sig_loopback =7319;
10075: waveform_sig_loopback =5734;
10076: waveform_sig_loopback =6769;
10077: waveform_sig_loopback =6629;
10078: waveform_sig_loopback =6774;
10079: waveform_sig_loopback =5751;
10080: waveform_sig_loopback =7885;
10081: waveform_sig_loopback =6169;
10082: waveform_sig_loopback =5821;
10083: waveform_sig_loopback =7962;
10084: waveform_sig_loopback =6276;
10085: waveform_sig_loopback =6109;
10086: waveform_sig_loopback =7347;
10087: waveform_sig_loopback =7151;
10088: waveform_sig_loopback =5835;
10089: waveform_sig_loopback =6890;
10090: waveform_sig_loopback =7825;
10091: waveform_sig_loopback =6214;
10092: waveform_sig_loopback =5809;
10093: waveform_sig_loopback =8163;
10094: waveform_sig_loopback =7352;
10095: waveform_sig_loopback =5068;
10096: waveform_sig_loopback =7540;
10097: waveform_sig_loopback =8286;
10098: waveform_sig_loopback =5174;
10099: waveform_sig_loopback =9200;
10100: waveform_sig_loopback =4930;
10101: waveform_sig_loopback =5171;
10102: waveform_sig_loopback =10342;
10103: waveform_sig_loopback =6319;
10104: waveform_sig_loopback =6278;
10105: waveform_sig_loopback =6190;
10106: waveform_sig_loopback =7276;
10107: waveform_sig_loopback =8960;
10108: waveform_sig_loopback =5815;
10109: waveform_sig_loopback =6181;
10110: waveform_sig_loopback =8283;
10111: waveform_sig_loopback =6215;
10112: waveform_sig_loopback =7955;
10113: waveform_sig_loopback =6187;
10114: waveform_sig_loopback =7179;
10115: waveform_sig_loopback =8129;
10116: waveform_sig_loopback =5946;
10117: waveform_sig_loopback =7527;
10118: waveform_sig_loopback =7238;
10119: waveform_sig_loopback =6986;
10120: waveform_sig_loopback =6567;
10121: waveform_sig_loopback =8322;
10122: waveform_sig_loopback =6416;
10123: waveform_sig_loopback =6647;
10124: waveform_sig_loopback =8197;
10125: waveform_sig_loopback =6682;
10126: waveform_sig_loopback =6746;
10127: waveform_sig_loopback =7596;
10128: waveform_sig_loopback =7647;
10129: waveform_sig_loopback =6259;
10130: waveform_sig_loopback =7148;
10131: waveform_sig_loopback =8431;
10132: waveform_sig_loopback =6404;
10133: waveform_sig_loopback =6101;
10134: waveform_sig_loopback =8897;
10135: waveform_sig_loopback =7286;
10136: waveform_sig_loopback =5481;
10137: waveform_sig_loopback =8268;
10138: waveform_sig_loopback =8050;
10139: waveform_sig_loopback =5896;
10140: waveform_sig_loopback =9441;
10141: waveform_sig_loopback =4723;
10142: waveform_sig_loopback =6232;
10143: waveform_sig_loopback =10160;
10144: waveform_sig_loopback =6584;
10145: waveform_sig_loopback =6796;
10146: waveform_sig_loopback =5914;
10147: waveform_sig_loopback =8111;
10148: waveform_sig_loopback =8955;
10149: waveform_sig_loopback =5726;
10150: waveform_sig_loopback =6924;
10151: waveform_sig_loopback =7985;
10152: waveform_sig_loopback =6640;
10153: waveform_sig_loopback =8243;
10154: waveform_sig_loopback =5874;
10155: waveform_sig_loopback =7776;
10156: waveform_sig_loopback =8031;
10157: waveform_sig_loopback =6017;
10158: waveform_sig_loopback =7849;
10159: waveform_sig_loopback =7169;
10160: waveform_sig_loopback =7105;
10161: waveform_sig_loopback =6759;
10162: waveform_sig_loopback =8287;
10163: waveform_sig_loopback =6352;
10164: waveform_sig_loopback =6977;
10165: waveform_sig_loopback =7985;
10166: waveform_sig_loopback =6831;
10167: waveform_sig_loopback =6805;
10168: waveform_sig_loopback =7347;
10169: waveform_sig_loopback =7966;
10170: waveform_sig_loopback =5920;
10171: waveform_sig_loopback =7144;
10172: waveform_sig_loopback =8701;
10173: waveform_sig_loopback =5807;
10174: waveform_sig_loopback =6403;
10175: waveform_sig_loopback =8794;
10176: waveform_sig_loopback =6757;
10177: waveform_sig_loopback =5852;
10178: waveform_sig_loopback =7819;
10179: waveform_sig_loopback =7808;
10180: waveform_sig_loopback =6072;
10181: waveform_sig_loopback =8858;
10182: waveform_sig_loopback =4692;
10183: waveform_sig_loopback =6147;
10184: waveform_sig_loopback =9636;
10185: waveform_sig_loopback =6706;
10186: waveform_sig_loopback =6138;
10187: waveform_sig_loopback =5807;
10188: waveform_sig_loopback =8046;
10189: waveform_sig_loopback =8254;
10190: waveform_sig_loopback =5622;
10191: waveform_sig_loopback =6665;
10192: waveform_sig_loopback =7456;
10193: waveform_sig_loopback =6413;
10194: waveform_sig_loopback =7591;
10195: waveform_sig_loopback =5628;
10196: waveform_sig_loopback =7659;
10197: waveform_sig_loopback =7199;
10198: waveform_sig_loopback =5595;
10199: waveform_sig_loopback =7680;
10200: waveform_sig_loopback =6592;
10201: waveform_sig_loopback =6632;
10202: waveform_sig_loopback =6319;
10203: waveform_sig_loopback =7724;
10204: waveform_sig_loopback =6102;
10205: waveform_sig_loopback =6329;
10206: waveform_sig_loopback =7271;
10207: waveform_sig_loopback =6686;
10208: waveform_sig_loopback =5920;
10209: waveform_sig_loopback =6966;
10210: waveform_sig_loopback =7492;
10211: waveform_sig_loopback =4950;
10212: waveform_sig_loopback =7177;
10213: waveform_sig_loopback =7690;
10214: waveform_sig_loopback =5023;
10215: waveform_sig_loopback =6420;
10216: waveform_sig_loopback =7598;
10217: waveform_sig_loopback =6378;
10218: waveform_sig_loopback =5218;
10219: waveform_sig_loopback =6967;
10220: waveform_sig_loopback =7568;
10221: waveform_sig_loopback =4935;
10222: waveform_sig_loopback =8350;
10223: waveform_sig_loopback =4024;
10224: waveform_sig_loopback =5270;
10225: waveform_sig_loopback =9198;
10226: waveform_sig_loopback =5704;
10227: waveform_sig_loopback =5305;
10228: waveform_sig_loopback =5398;
10229: waveform_sig_loopback =7086;
10230: waveform_sig_loopback =7506;
10231: waveform_sig_loopback =4841;
10232: waveform_sig_loopback =5922;
10233: waveform_sig_loopback =6588;
10234: waveform_sig_loopback =5827;
10235: waveform_sig_loopback =6695;
10236: waveform_sig_loopback =4701;
10237: waveform_sig_loopback =7031;
10238: waveform_sig_loopback =5989;
10239: waveform_sig_loopback =5203;
10240: waveform_sig_loopback =6583;
10241: waveform_sig_loopback =5393;
10242: waveform_sig_loopback =6281;
10243: waveform_sig_loopback =5062;
10244: waveform_sig_loopback =6875;
10245: waveform_sig_loopback =5243;
10246: waveform_sig_loopback =5031;
10247: waveform_sig_loopback =6882;
10248: waveform_sig_loopback =5274;
10249: waveform_sig_loopback =4894;
10250: waveform_sig_loopback =6543;
10251: waveform_sig_loopback =5799;
10252: waveform_sig_loopback =4302;
10253: waveform_sig_loopback =6197;
10254: waveform_sig_loopback =6348;
10255: waveform_sig_loopback =4322;
10256: waveform_sig_loopback =5097;
10257: waveform_sig_loopback =6640;
10258: waveform_sig_loopback =5394;
10259: waveform_sig_loopback =3918;
10260: waveform_sig_loopback =6094;
10261: waveform_sig_loopback =6335;
10262: waveform_sig_loopback =3790;
10263: waveform_sig_loopback =7376;
10264: waveform_sig_loopback =2611;
10265: waveform_sig_loopback =4356;
10266: waveform_sig_loopback =8145;
10267: waveform_sig_loopback =4381;
10268: waveform_sig_loopback =4083;
10269: waveform_sig_loopback =4419;
10270: waveform_sig_loopback =5818;
10271: waveform_sig_loopback =6241;
10272: waveform_sig_loopback =3761;
10273: waveform_sig_loopback =4493;
10274: waveform_sig_loopback =5604;
10275: waveform_sig_loopback =4562;
10276: waveform_sig_loopback =5152;
10277: waveform_sig_loopback =3896;
10278: waveform_sig_loopback =5487;
10279: waveform_sig_loopback =4733;
10280: waveform_sig_loopback =4186;
10281: waveform_sig_loopback =4794;
10282: waveform_sig_loopback =4578;
10283: waveform_sig_loopback =4695;
10284: waveform_sig_loopback =3626;
10285: waveform_sig_loopback =6056;
10286: waveform_sig_loopback =3296;
10287: waveform_sig_loopback =4098;
10288: waveform_sig_loopback =5579;
10289: waveform_sig_loopback =3526;
10290: waveform_sig_loopback =3957;
10291: waveform_sig_loopback =4949;
10292: waveform_sig_loopback =4401;
10293: waveform_sig_loopback =3103;
10294: waveform_sig_loopback =4623;
10295: waveform_sig_loopback =5041;
10296: waveform_sig_loopback =2882;
10297: waveform_sig_loopback =3629;
10298: waveform_sig_loopback =5338;
10299: waveform_sig_loopback =3895;
10300: waveform_sig_loopback =2316;
10301: waveform_sig_loopback =4927;
10302: waveform_sig_loopback =4671;
10303: waveform_sig_loopback =2296;
10304: waveform_sig_loopback =6117;
10305: waveform_sig_loopback =721;
10306: waveform_sig_loopback =3211;
10307: waveform_sig_loopback =6733;
10308: waveform_sig_loopback =2486;
10309: waveform_sig_loopback =2835;
10310: waveform_sig_loopback =2882;
10311: waveform_sig_loopback =4124;
10312: waveform_sig_loopback =5055;
10313: waveform_sig_loopback =1762;
10314: waveform_sig_loopback =3085;
10315: waveform_sig_loopback =4254;
10316: waveform_sig_loopback =2566;
10317: waveform_sig_loopback =3955;
10318: waveform_sig_loopback =2138;
10319: waveform_sig_loopback =3717;
10320: waveform_sig_loopback =3572;
10321: waveform_sig_loopback =2169;
10322: waveform_sig_loopback =3368;
10323: waveform_sig_loopback =3173;
10324: waveform_sig_loopback =2621;
10325: waveform_sig_loopback =2521;
10326: waveform_sig_loopback =4141;
10327: waveform_sig_loopback =1555;
10328: waveform_sig_loopback =2814;
10329: waveform_sig_loopback =3555;
10330: waveform_sig_loopback =2053;
10331: waveform_sig_loopback =2280;
10332: waveform_sig_loopback =3242;
10333: waveform_sig_loopback =2703;
10334: waveform_sig_loopback =1465;
10335: waveform_sig_loopback =2933;
10336: waveform_sig_loopback =3317;
10337: waveform_sig_loopback =1247;
10338: waveform_sig_loopback =1704;
10339: waveform_sig_loopback =3999;
10340: waveform_sig_loopback =1874;
10341: waveform_sig_loopback =539;
10342: waveform_sig_loopback =3728;
10343: waveform_sig_loopback =2289;
10344: waveform_sig_loopback =1053;
10345: waveform_sig_loopback =4316;
10346: waveform_sig_loopback =-1546;
10347: waveform_sig_loopback =2331;
10348: waveform_sig_loopback =4354;
10349: waveform_sig_loopback =778;
10350: waveform_sig_loopback =1374;
10351: waveform_sig_loopback =607;
10352: waveform_sig_loopback =2904;
10353: waveform_sig_loopback =2993;
10354: waveform_sig_loopback =-286;
10355: waveform_sig_loopback =1875;
10356: waveform_sig_loopback =1957;
10357: waveform_sig_loopback =1019;
10358: waveform_sig_loopback =2265;
10359: waveform_sig_loopback =-19;
10360: waveform_sig_loopback =2354;
10361: waveform_sig_loopback =1486;
10362: waveform_sig_loopback =316;
10363: waveform_sig_loopback =1776;
10364: waveform_sig_loopback =1178;
10365: waveform_sig_loopback =756;
10366: waveform_sig_loopback =865;
10367: waveform_sig_loopback =2120;
10368: waveform_sig_loopback =-334;
10369: waveform_sig_loopback =1263;
10370: waveform_sig_loopback =1369;
10371: waveform_sig_loopback =365;
10372: waveform_sig_loopback =500;
10373: waveform_sig_loopback =1128;
10374: waveform_sig_loopback =1187;
10375: waveform_sig_loopback =-728;
10376: waveform_sig_loopback =1165;
10377: waveform_sig_loopback =1688;
10378: waveform_sig_loopback =-1087;
10379: waveform_sig_loopback =303;
10380: waveform_sig_loopback =2009;
10381: waveform_sig_loopback =-321;
10382: waveform_sig_loopback =-899;
10383: waveform_sig_loopback =1621;
10384: waveform_sig_loopback =282;
10385: waveform_sig_loopback =-417;
10386: waveform_sig_loopback =1991;
10387: waveform_sig_loopback =-3266;
10388: waveform_sig_loopback =703;
10389: waveform_sig_loopback =2096;
10390: waveform_sig_loopback =-713;
10391: waveform_sig_loopback =-822;
10392: waveform_sig_loopback =-1213;
10393: waveform_sig_loopback =1380;
10394: waveform_sig_loopback =693;
10395: waveform_sig_loopback =-2011;
10396: waveform_sig_loopback =68;
10397: waveform_sig_loopback =-225;
10398: waveform_sig_loopback =-521;
10399: waveform_sig_loopback =177;
10400: waveform_sig_loopback =-2001;
10401: waveform_sig_loopback =798;
10402: waveform_sig_loopback =-746;
10403: waveform_sig_loopback =-1447;
10404: waveform_sig_loopback =6;
10405: waveform_sig_loopback =-998;
10406: waveform_sig_loopback =-912;
10407: waveform_sig_loopback =-944;
10408: waveform_sig_loopback =-90;
10409: waveform_sig_loopback =-1936;
10410: waveform_sig_loopback =-730;
10411: waveform_sig_loopback =-567;
10412: waveform_sig_loopback =-1203;
10413: waveform_sig_loopback =-1798;
10414: waveform_sig_loopback =-368;
10415: waveform_sig_loopback =-814;
10416: waveform_sig_loopback =-2908;
10417: waveform_sig_loopback =-186;
10418: waveform_sig_loopback =-577;
10419: waveform_sig_loopback =-2962;
10420: waveform_sig_loopback =-1217;
10421: waveform_sig_loopback =-269;
10422: waveform_sig_loopback =-2019;
10423: waveform_sig_loopback =-2744;
10424: waveform_sig_loopback =-404;
10425: waveform_sig_loopback =-1431;
10426: waveform_sig_loopback =-2350;
10427: waveform_sig_loopback =-23;
10428: waveform_sig_loopback =-5068;
10429: waveform_sig_loopback =-1139;
10430: waveform_sig_loopback =163;
10431: waveform_sig_loopback =-2548;
10432: waveform_sig_loopback =-2977;
10433: waveform_sig_loopback =-2760;
10434: waveform_sig_loopback =-471;
10435: waveform_sig_loopback =-1533;
10436: waveform_sig_loopback =-3562;
10437: waveform_sig_loopback =-1907;
10438: waveform_sig_loopback =-2136;
10439: waveform_sig_loopback =-2161;
10440: waveform_sig_loopback =-2095;
10441: waveform_sig_loopback =-3505;
10442: waveform_sig_loopback =-989;
10443: waveform_sig_loopback =-2967;
10444: waveform_sig_loopback =-2888;
10445: waveform_sig_loopback =-2015;
10446: waveform_sig_loopback =-2877;
10447: waveform_sig_loopback =-2550;
10448: waveform_sig_loopback =-3063;
10449: waveform_sig_loopback =-1710;
10450: waveform_sig_loopback =-3707;
10451: waveform_sig_loopback =-2842;
10452: waveform_sig_loopback =-2024;
10453: waveform_sig_loopback =-3310;
10454: waveform_sig_loopback =-3594;
10455: waveform_sig_loopback =-1869;
10456: waveform_sig_loopback =-3090;
10457: waveform_sig_loopback =-4351;
10458: waveform_sig_loopback =-1966;
10459: waveform_sig_loopback =-2741;
10460: waveform_sig_loopback =-4544;
10461: waveform_sig_loopback =-3028;
10462: waveform_sig_loopback =-2113;
10463: waveform_sig_loopback =-3770;
10464: waveform_sig_loopback =-4576;
10465: waveform_sig_loopback =-2101;
10466: waveform_sig_loopback =-3208;
10467: waveform_sig_loopback =-4217;
10468: waveform_sig_loopback =-1797;
10469: waveform_sig_loopback =-6788;
10470: waveform_sig_loopback =-2945;
10471: waveform_sig_loopback =-1373;
10472: waveform_sig_loopback =-4482;
10473: waveform_sig_loopback =-4886;
10474: waveform_sig_loopback =-4084;
10475: waveform_sig_loopback =-2606;
10476: waveform_sig_loopback =-3068;
10477: waveform_sig_loopback =-5177;
10478: waveform_sig_loopback =-3935;
10479: waveform_sig_loopback =-3475;
10480: waveform_sig_loopback =-4083;
10481: waveform_sig_loopback =-3871;
10482: waveform_sig_loopback =-4899;
10483: waveform_sig_loopback =-3058;
10484: waveform_sig_loopback =-4448;
10485: waveform_sig_loopback =-4420;
10486: waveform_sig_loopback =-3994;
10487: waveform_sig_loopback =-4164;
10488: waveform_sig_loopback =-4481;
10489: waveform_sig_loopback =-4629;
10490: waveform_sig_loopback =-3201;
10491: waveform_sig_loopback =-5542;
10492: waveform_sig_loopback =-4285;
10493: waveform_sig_loopback =-3599;
10494: waveform_sig_loopback =-5134;
10495: waveform_sig_loopback =-5025;
10496: waveform_sig_loopback =-3319;
10497: waveform_sig_loopback =-5032;
10498: waveform_sig_loopback =-5585;
10499: waveform_sig_loopback =-3612;
10500: waveform_sig_loopback =-4441;
10501: waveform_sig_loopback =-5755;
10502: waveform_sig_loopback =-4911;
10503: waveform_sig_loopback =-3441;
10504: waveform_sig_loopback =-5344;
10505: waveform_sig_loopback =-6337;
10506: waveform_sig_loopback =-3123;
10507: waveform_sig_loopback =-5124;
10508: waveform_sig_loopback =-5580;
10509: waveform_sig_loopback =-3165;
10510: waveform_sig_loopback =-8718;
10511: waveform_sig_loopback =-3951;
10512: waveform_sig_loopback =-2932;
10513: waveform_sig_loopback =-6278;
10514: waveform_sig_loopback =-5996;
10515: waveform_sig_loopback =-5624;
10516: waveform_sig_loopback =-4083;
10517: waveform_sig_loopback =-4313;
10518: waveform_sig_loopback =-6995;
10519: waveform_sig_loopback =-5051;
10520: waveform_sig_loopback =-4876;
10521: waveform_sig_loopback =-5682;
10522: waveform_sig_loopback =-5012;
10523: waveform_sig_loopback =-6407;
10524: waveform_sig_loopback =-4457;
10525: waveform_sig_loopback =-5634;
10526: waveform_sig_loopback =-6010;
10527: waveform_sig_loopback =-5307;
10528: waveform_sig_loopback =-5359;
10529: waveform_sig_loopback =-6104;
10530: waveform_sig_loopback =-5741;
10531: waveform_sig_loopback =-4559;
10532: waveform_sig_loopback =-7176;
10533: waveform_sig_loopback =-5296;
10534: waveform_sig_loopback =-5138;
10535: waveform_sig_loopback =-6532;
10536: waveform_sig_loopback =-6043;
10537: waveform_sig_loopback =-4948;
10538: waveform_sig_loopback =-6191;
10539: waveform_sig_loopback =-6780;
10540: waveform_sig_loopback =-5127;
10541: waveform_sig_loopback =-5489;
10542: waveform_sig_loopback =-7161;
10543: waveform_sig_loopback =-6289;
10544: waveform_sig_loopback =-4463;
10545: waveform_sig_loopback =-6825;
10546: waveform_sig_loopback =-7346;
10547: waveform_sig_loopback =-4279;
10548: waveform_sig_loopback =-6952;
10549: waveform_sig_loopback =-6038;
10550: waveform_sig_loopback =-4560;
10551: waveform_sig_loopback =-10163;
10552: waveform_sig_loopback =-4660;
10553: waveform_sig_loopback =-4380;
10554: waveform_sig_loopback =-7264;
10555: waveform_sig_loopback =-7138;
10556: waveform_sig_loopback =-7021;
10557: waveform_sig_loopback =-4796;
10558: waveform_sig_loopback =-5525;
10559: waveform_sig_loopback =-8410;
10560: waveform_sig_loopback =-5700;
10561: waveform_sig_loopback =-6255;
10562: waveform_sig_loopback =-6632;
10563: waveform_sig_loopback =-6000;
10564: waveform_sig_loopback =-7811;
10565: waveform_sig_loopback =-5119;
10566: waveform_sig_loopback =-6853;
10567: waveform_sig_loopback =-7177;
10568: waveform_sig_loopback =-6093;
10569: waveform_sig_loopback =-6453;
10570: waveform_sig_loopback =-7194;
10571: waveform_sig_loopback =-6514;
10572: waveform_sig_loopback =-5757;
10573: waveform_sig_loopback =-8020;
10574: waveform_sig_loopback =-5984;
10575: waveform_sig_loopback =-6557;
10576: waveform_sig_loopback =-7101;
10577: waveform_sig_loopback =-6962;
10578: waveform_sig_loopback =-6104;
10579: waveform_sig_loopback =-6758;
10580: waveform_sig_loopback =-7988;
10581: waveform_sig_loopback =-5747;
10582: waveform_sig_loopback =-6292;
10583: waveform_sig_loopback =-8384;
10584: waveform_sig_loopback =-6529;
10585: waveform_sig_loopback =-5474;
10586: waveform_sig_loopback =-7942;
10587: waveform_sig_loopback =-7814;
10588: waveform_sig_loopback =-5178;
10589: waveform_sig_loopback =-7597;
10590: waveform_sig_loopback =-6747;
10591: waveform_sig_loopback =-5774;
10592: waveform_sig_loopback =-10636;
10593: waveform_sig_loopback =-5044;
10594: waveform_sig_loopback =-5651;
10595: waveform_sig_loopback =-7854;
10596: waveform_sig_loopback =-7811;
10597: waveform_sig_loopback =-7772;
10598: waveform_sig_loopback =-5163;
10599: waveform_sig_loopback =-6667;
10600: waveform_sig_loopback =-8827;
10601: waveform_sig_loopback =-6098;
10602: waveform_sig_loopback =-7411;
10603: waveform_sig_loopback =-6747;
10604: waveform_sig_loopback =-6901;
10605: waveform_sig_loopback =-8394;
10606: waveform_sig_loopback =-5416;
10607: waveform_sig_loopback =-7925;
10608: waveform_sig_loopback =-7317;
10609: waveform_sig_loopback =-6714;
10610: waveform_sig_loopback =-7254;
10611: waveform_sig_loopback =-7420;
10612: waveform_sig_loopback =-7089;
10613: waveform_sig_loopback =-6356;
10614: waveform_sig_loopback =-8420;
10615: waveform_sig_loopback =-6543;
10616: waveform_sig_loopback =-6901;
10617: waveform_sig_loopback =-7575;
10618: waveform_sig_loopback =-7550;
10619: waveform_sig_loopback =-6404;
10620: waveform_sig_loopback =-7198;
10621: waveform_sig_loopback =-8541;
10622: waveform_sig_loopback =-5947;
10623: waveform_sig_loopback =-6838;
10624: waveform_sig_loopback =-8925;
10625: waveform_sig_loopback =-6483;
10626: waveform_sig_loopback =-6209;
10627: waveform_sig_loopback =-8183;
10628: waveform_sig_loopback =-7903;
10629: waveform_sig_loopback =-5856;
10630: waveform_sig_loopback =-7659;
10631: waveform_sig_loopback =-7076;
10632: waveform_sig_loopback =-6279;
10633: waveform_sig_loopback =-10583;
10634: waveform_sig_loopback =-5508;
10635: waveform_sig_loopback =-5748;
10636: waveform_sig_loopback =-7989;
10637: waveform_sig_loopback =-8386;
10638: waveform_sig_loopback =-7552;
10639: waveform_sig_loopback =-5523;
10640: waveform_sig_loopback =-7024;
10641: waveform_sig_loopback =-8689;
10642: waveform_sig_loopback =-6562;
10643: waveform_sig_loopback =-7436;
10644: waveform_sig_loopback =-6783;
10645: waveform_sig_loopback =-7351;
10646: waveform_sig_loopback =-8195;
10647: waveform_sig_loopback =-5632;
10648: waveform_sig_loopback =-8131;
10649: waveform_sig_loopback =-7144;
10650: waveform_sig_loopback =-6990;
10651: waveform_sig_loopback =-7249;
10652: waveform_sig_loopback =-7420;
10653: waveform_sig_loopback =-7158;
10654: waveform_sig_loopback =-6439;
10655: waveform_sig_loopback =-8284;
10656: waveform_sig_loopback =-6695;
10657: waveform_sig_loopback =-6788;
10658: waveform_sig_loopback =-7522;
10659: waveform_sig_loopback =-7679;
10660: waveform_sig_loopback =-5920;
10661: waveform_sig_loopback =-7551;
10662: waveform_sig_loopback =-8284;
10663: waveform_sig_loopback =-5507;
10664: waveform_sig_loopback =-7267;
10665: waveform_sig_loopback =-8357;
10666: waveform_sig_loopback =-6420;
10667: waveform_sig_loopback =-6258;
10668: waveform_sig_loopback =-7698;
10669: waveform_sig_loopback =-8080;
10670: waveform_sig_loopback =-5401;
10671: waveform_sig_loopback =-7493;
10672: waveform_sig_loopback =-7041;
10673: waveform_sig_loopback =-5915;
10674: waveform_sig_loopback =-10539;
10675: waveform_sig_loopback =-5070;
10676: waveform_sig_loopback =-5424;
10677: waveform_sig_loopback =-8142;
10678: waveform_sig_loopback =-7893;
10679: waveform_sig_loopback =-7082;
10680: waveform_sig_loopback =-5497;
10681: waveform_sig_loopback =-6610;
10682: waveform_sig_loopback =-8433;
10683: waveform_sig_loopback =-6206;
10684: waveform_sig_loopback =-6993;
10685: waveform_sig_loopback =-6584;
10686: waveform_sig_loopback =-6984;
10687: waveform_sig_loopback =-7566;
10688: waveform_sig_loopback =-5468;
10689: waveform_sig_loopback =-7691;
10690: waveform_sig_loopback =-6649;
10691: waveform_sig_loopback =-6686;
10692: waveform_sig_loopback =-6710;
10693: waveform_sig_loopback =-6994;
10694: waveform_sig_loopback =-6805;
10695: waveform_sig_loopback =-5764;
10696: waveform_sig_loopback =-7977;
10697: waveform_sig_loopback =-6258;
10698: waveform_sig_loopback =-5921;
10699: waveform_sig_loopback =-7555;
10700: waveform_sig_loopback =-6695;
10701: waveform_sig_loopback =-5479;
10702: waveform_sig_loopback =-7415;
10703: waveform_sig_loopback =-7062;
10704: waveform_sig_loopback =-5510;
10705: waveform_sig_loopback =-6539;
10706: waveform_sig_loopback =-7570;
10707: waveform_sig_loopback =-6142;
10708: waveform_sig_loopback =-5273;
10709: waveform_sig_loopback =-7424;
10710: waveform_sig_loopback =-7320;
10711: waveform_sig_loopback =-4450;
10712: waveform_sig_loopback =-7342;
10713: waveform_sig_loopback =-5896;
10714: waveform_sig_loopback =-5436;
10715: waveform_sig_loopback =-9971;
10716: waveform_sig_loopback =-3958;
10717: waveform_sig_loopback =-4995;
10718: waveform_sig_loopback =-7397;
10719: waveform_sig_loopback =-7070;
10720: waveform_sig_loopback =-6323;
10721: waveform_sig_loopback =-4708;
10722: waveform_sig_loopback =-5878;
10723: waveform_sig_loopback =-7669;
10724: waveform_sig_loopback =-5416;
10725: waveform_sig_loopback =-6018;
10726: waveform_sig_loopback =-5918;
10727: waveform_sig_loopback =-6175;
10728: waveform_sig_loopback =-6509;
10729: waveform_sig_loopback =-4944;
10730: waveform_sig_loopback =-6525;
10731: waveform_sig_loopback =-5907;
10732: waveform_sig_loopback =-5972;
10733: waveform_sig_loopback =-5338;
10734: waveform_sig_loopback =-6672;
10735: waveform_sig_loopback =-5461;
10736: waveform_sig_loopback =-4881;
10737: waveform_sig_loopback =-7431;
10738: waveform_sig_loopback =-4594;
10739: waveform_sig_loopback =-5564;
10740: waveform_sig_loopback =-6371;
10741: waveform_sig_loopback =-5478;
10742: waveform_sig_loopback =-4970;
10743: waveform_sig_loopback =-5978;
10744: waveform_sig_loopback =-6280;
10745: waveform_sig_loopback =-4382;
10746: waveform_sig_loopback =-5435;
10747: waveform_sig_loopback =-6808;
10748: waveform_sig_loopback =-4756;
10749: waveform_sig_loopback =-4345;
10750: waveform_sig_loopback =-6430;
10751: waveform_sig_loopback =-6133;
10752: waveform_sig_loopback =-3310;
10753: waveform_sig_loopback =-6376;
10754: waveform_sig_loopback =-4673;
10755: waveform_sig_loopback =-4399;
10756: waveform_sig_loopback =-8944;
10757: waveform_sig_loopback =-2470;
10758: waveform_sig_loopback =-4062;
10759: waveform_sig_loopback =-6352;
10760: waveform_sig_loopback =-5587;
10761: waveform_sig_loopback =-5401;
10762: waveform_sig_loopback =-3321;
10763: waveform_sig_loopback =-4637;
10764: waveform_sig_loopback =-6774;
10765: waveform_sig_loopback =-3716;
10766: waveform_sig_loopback =-5111;
10767: waveform_sig_loopback =-4682;
10768: waveform_sig_loopback =-4657;
10769: waveform_sig_loopback =-5644;
10770: waveform_sig_loopback =-3402;
10771: waveform_sig_loopback =-5299;
10772: waveform_sig_loopback =-4893;
10773: waveform_sig_loopback =-4243;
10774: waveform_sig_loopback =-4361;
10775: waveform_sig_loopback =-5332;
10776: waveform_sig_loopback =-3779;
10777: waveform_sig_loopback =-4070;
10778: waveform_sig_loopback =-5716;
10779: waveform_sig_loopback =-3323;
10780: waveform_sig_loopback =-4388;
10781: waveform_sig_loopback =-4784;
10782: waveform_sig_loopback =-4271;
10783: waveform_sig_loopback =-3469;
10784: waveform_sig_loopback =-4662;
10785: waveform_sig_loopback =-4911;
10786: waveform_sig_loopback =-2865;
10787: waveform_sig_loopback =-4099;
10788: waveform_sig_loopback =-5444;
10789: waveform_sig_loopback =-3227;
10790: waveform_sig_loopback =-2824;
10791: waveform_sig_loopback =-5253;
10792: waveform_sig_loopback =-4441;
10793: waveform_sig_loopback =-1813;
10794: waveform_sig_loopback =-5223;
10795: waveform_sig_loopback =-2702;
10796: waveform_sig_loopback =-3453;
10797: waveform_sig_loopback =-7278;
10798: waveform_sig_loopback =-557;
10799: waveform_sig_loopback =-3216;
10800: waveform_sig_loopback =-4397;
10801: waveform_sig_loopback =-4209;
10802: waveform_sig_loopback =-4034;
10803: waveform_sig_loopback =-1304;
10804: waveform_sig_loopback =-3714;
10805: waveform_sig_loopback =-4901;
10806: waveform_sig_loopback =-2029;
10807: waveform_sig_loopback =-3981;
10808: waveform_sig_loopback =-2615;
10809: waveform_sig_loopback =-3434;
10810: waveform_sig_loopback =-3969;
10811: waveform_sig_loopback =-1548;
10812: waveform_sig_loopback =-4141;
10813: waveform_sig_loopback =-2964;
10814: waveform_sig_loopback =-2653;
10815: waveform_sig_loopback =-2989;
10816: waveform_sig_loopback =-3448;
10817: waveform_sig_loopback =-2224;
10818: waveform_sig_loopback =-2584;
10819: waveform_sig_loopback =-3898;
10820: waveform_sig_loopback =-1750;
10821: waveform_sig_loopback =-2766;
10822: waveform_sig_loopback =-3073;
10823: waveform_sig_loopback =-2658;
10824: waveform_sig_loopback =-1743;
10825: waveform_sig_loopback =-2930;
10826: waveform_sig_loopback =-3356;
10827: waveform_sig_loopback =-988;
10828: waveform_sig_loopback =-2452;
10829: waveform_sig_loopback =-3986;
10830: waveform_sig_loopback =-1033;
10831: waveform_sig_loopback =-1441;
10832: waveform_sig_loopback =-3646;
10833: waveform_sig_loopback =-2267;
10834: waveform_sig_loopback =-597;
10835: waveform_sig_loopback =-3165;
10836: waveform_sig_loopback =-826;
10837: waveform_sig_loopback =-2298;
10838: waveform_sig_loopback =-4821;
10839: waveform_sig_loopback =821;
10840: waveform_sig_loopback =-1365;
10841: waveform_sig_loopback =-2408;
10842: waveform_sig_loopback =-2976;
10843: waveform_sig_loopback =-1684;
10844: waveform_sig_loopback =364;
10845: waveform_sig_loopback =-2222;
10846: waveform_sig_loopback =-2710;
10847: waveform_sig_loopback =-568;
10848: waveform_sig_loopback =-2025;
10849: waveform_sig_loopback =-621;
10850: waveform_sig_loopback =-2031;
10851: waveform_sig_loopback =-1746;
10852: waveform_sig_loopback =179;
10853: waveform_sig_loopback =-2450;
10854: waveform_sig_loopback =-865;
10855: waveform_sig_loopback =-978;
10856: waveform_sig_loopback =-1172;
10857: waveform_sig_loopback =-1489;
10858: waveform_sig_loopback =-390;
10859: waveform_sig_loopback =-905;
10860: waveform_sig_loopback =-1755;
10861: waveform_sig_loopback =-189;
10862: waveform_sig_loopback =-699;
10863: waveform_sig_loopback =-1227;
10864: waveform_sig_loopback =-1060;
10865: waveform_sig_loopback =589;
10866: waveform_sig_loopback =-1594;
10867: waveform_sig_loopback =-1309;
10868: waveform_sig_loopback =1062;
10869: waveform_sig_loopback =-1083;
10870: waveform_sig_loopback =-1679;
10871: waveform_sig_loopback =659;
10872: waveform_sig_loopback =277;
10873: waveform_sig_loopback =-1542;
10874: waveform_sig_loopback =-528;
10875: waveform_sig_loopback =1299;
10876: waveform_sig_loopback =-1231;
10877: waveform_sig_loopback =948;
10878: waveform_sig_loopback =-519;
10879: waveform_sig_loopback =-2737;
10880: waveform_sig_loopback =2517;
10881: waveform_sig_loopback =644;
10882: waveform_sig_loopback =-723;
10883: waveform_sig_loopback =-1149;
10884: waveform_sig_loopback =599;
10885: waveform_sig_loopback =1776;
10886: waveform_sig_loopback =-115;
10887: waveform_sig_loopback =-758;
10888: waveform_sig_loopback =1028;
10889: waveform_sig_loopback =179;
10890: waveform_sig_loopback =1034;
10891: waveform_sig_loopback =-197;
10892: waveform_sig_loopback =193;
10893: waveform_sig_loopback =1820;
10894: waveform_sig_loopback =-351;
10895: waveform_sig_loopback =1091;
10896: waveform_sig_loopback =493;
10897: waveform_sig_loopback =845;
10898: waveform_sig_loopback =622;
10899: waveform_sig_loopback =1304;
10900: waveform_sig_loopback =1024;
10901: waveform_sig_loopback =-29;
10902: waveform_sig_loopback =1863;
10903: waveform_sig_loopback =1390;
10904: waveform_sig_loopback =155;
10905: waveform_sig_loopback =1190;
10906: waveform_sig_loopback =2515;
10907: waveform_sig_loopback =-41;
10908: waveform_sig_loopback =1003;
10909: waveform_sig_loopback =2726;
10910: waveform_sig_loopback =781;
10911: waveform_sig_loopback =461;
10912: waveform_sig_loopback =2275;
10913: waveform_sig_loopback =2294;
10914: waveform_sig_loopback =405;
10915: waveform_sig_loopback =1161;
10916: waveform_sig_loopback =3423;
10917: waveform_sig_loopback =476;
10918: waveform_sig_loopback =2932;
10919: waveform_sig_loopback =1421;
10920: waveform_sig_loopback =-1044;
10921: waveform_sig_loopback =4682;
10922: waveform_sig_loopback =2530;
10923: waveform_sig_loopback =784;
10924: waveform_sig_loopback =1037;
10925: waveform_sig_loopback =2434;
10926: waveform_sig_loopback =3485;
10927: waveform_sig_loopback =1906;
10928: waveform_sig_loopback =869;
10929: waveform_sig_loopback =3074;
10930: waveform_sig_loopback =2116;
10931: waveform_sig_loopback =2617;
10932: waveform_sig_loopback =1817;
10933: waveform_sig_loopback =2293;
10934: waveform_sig_loopback =3369;
10935: waveform_sig_loopback =1595;
10936: waveform_sig_loopback =2820;
10937: waveform_sig_loopback =2462;
10938: waveform_sig_loopback =2891;
10939: waveform_sig_loopback =1910;
10940: waveform_sig_loopback =3432;
10941: waveform_sig_loopback =2950;
10942: waveform_sig_loopback =1563;
10943: waveform_sig_loopback =3847;
10944: waveform_sig_loopback =3009;
10945: waveform_sig_loopback =1984;
10946: waveform_sig_loopback =3306;
10947: waveform_sig_loopback =3870;
10948: waveform_sig_loopback =1815;
10949: waveform_sig_loopback =3087;
10950: waveform_sig_loopback =4140;
10951: waveform_sig_loopback =2651;
10952: waveform_sig_loopback =2260;
10953: waveform_sig_loopback =3990;
10954: waveform_sig_loopback =4228;
10955: waveform_sig_loopback =1792;
10956: waveform_sig_loopback =3134;
10957: waveform_sig_loopback =5422;
10958: waveform_sig_loopback =1680;
10959: waveform_sig_loopback =5118;
10960: waveform_sig_loopback =2866;
10961: waveform_sig_loopback =691;
10962: waveform_sig_loopback =6839;
10963: waveform_sig_loopback =3760;
10964: waveform_sig_loopback =2655;
10965: waveform_sig_loopback =2978;
10966: waveform_sig_loopback =3860;
10967: waveform_sig_loopback =5501;
10968: waveform_sig_loopback =3397;
10969: waveform_sig_loopback =2493;
10970: waveform_sig_loopback =5058;
10971: waveform_sig_loopback =3563;
10972: waveform_sig_loopback =4394;
10973: waveform_sig_loopback =3556;
10974: waveform_sig_loopback =3842;
10975: waveform_sig_loopback =5108;
10976: waveform_sig_loopback =3306;
10977: waveform_sig_loopback =4329;
10978: waveform_sig_loopback =4274;
10979: waveform_sig_loopback =4527;
10980: waveform_sig_loopback =3366;
10981: waveform_sig_loopback =5391;
10982: waveform_sig_loopback =4277;
10983: waveform_sig_loopback =3203;
10984: waveform_sig_loopback =5775;
10985: waveform_sig_loopback =4147;
10986: waveform_sig_loopback =3869;
10987: waveform_sig_loopback =4976;
10988: waveform_sig_loopback =5120;
10989: waveform_sig_loopback =3834;
10990: waveform_sig_loopback =4392;
10991: waveform_sig_loopback =5845;
10992: waveform_sig_loopback =4410;
10993: waveform_sig_loopback =3410;
10994: waveform_sig_loopback =6054;
10995: waveform_sig_loopback =5597;
10996: waveform_sig_loopback =3108;
10997: waveform_sig_loopback =5245;
10998: waveform_sig_loopback =6483;
10999: waveform_sig_loopback =3311;
11000: waveform_sig_loopback =6868;
11001: waveform_sig_loopback =3839;
11002: waveform_sig_loopback =2599;
11003: waveform_sig_loopback =8283;
11004: waveform_sig_loopback =4983;
11005: waveform_sig_loopback =4365;
11006: waveform_sig_loopback =4289;
11007: waveform_sig_loopback =5322;
11008: waveform_sig_loopback =7191;
11009: waveform_sig_loopback =4537;
11010: waveform_sig_loopback =4069;
11011: waveform_sig_loopback =6620;
11012: waveform_sig_loopback =4653;
11013: waveform_sig_loopback =6150;
11014: waveform_sig_loopback =4818;
11015: waveform_sig_loopback =5161;
11016: waveform_sig_loopback =6788;
11017: waveform_sig_loopback =4437;
11018: waveform_sig_loopback =5762;
11019: waveform_sig_loopback =5836;
11020: waveform_sig_loopback =5540;
11021: waveform_sig_loopback =4971;
11022: waveform_sig_loopback =6846;
11023: waveform_sig_loopback =5134;
11024: waveform_sig_loopback =5095;
11025: waveform_sig_loopback =6797;
11026: waveform_sig_loopback =5391;
11027: waveform_sig_loopback =5479;
11028: waveform_sig_loopback =5897;
11029: waveform_sig_loopback =6718;
11030: waveform_sig_loopback =4962;
11031: waveform_sig_loopback =5535;
11032: waveform_sig_loopback =7418;
11033: waveform_sig_loopback =5292;
11034: waveform_sig_loopback =4791;
11035: waveform_sig_loopback =7461;
11036: waveform_sig_loopback =6496;
11037: waveform_sig_loopback =4431;
11038: waveform_sig_loopback =6584;
11039: waveform_sig_loopback =7375;
11040: waveform_sig_loopback =4712;
11041: waveform_sig_loopback =8122;
11042: waveform_sig_loopback =4605;
11043: waveform_sig_loopback =4259;
11044: waveform_sig_loopback =9252;
11045: waveform_sig_loopback =6017;
11046: waveform_sig_loopback =5715;
11047: waveform_sig_loopback =5126;
11048: waveform_sig_loopback =6710;
11049: waveform_sig_loopback =8275;
11050: waveform_sig_loopback =5237;
11051: waveform_sig_loopback =5619;
11052: waveform_sig_loopback =7481;
11053: waveform_sig_loopback =5606;
11054: waveform_sig_loopback =7528;
11055: waveform_sig_loopback =5360;
11056: waveform_sig_loopback =6589;
11057: waveform_sig_loopback =7744;
11058: waveform_sig_loopback =5074;
11059: waveform_sig_loopback =7263;
11060: waveform_sig_loopback =6518;
11061: waveform_sig_loopback =6493;
11062: waveform_sig_loopback =6251;
11063: waveform_sig_loopback =7437;
11064: waveform_sig_loopback =6275;
11065: waveform_sig_loopback =6082;
11066: waveform_sig_loopback =7525;
11067: waveform_sig_loopback =6619;
11068: waveform_sig_loopback =6175;
11069: waveform_sig_loopback =6861;
11070: waveform_sig_loopback =7762;
11071: waveform_sig_loopback =5588;
11072: waveform_sig_loopback =6597;
11073: waveform_sig_loopback =8334;
11074: waveform_sig_loopback =5863;
11075: waveform_sig_loopback =5859;
11076: waveform_sig_loopback =8321;
11077: waveform_sig_loopback =7039;
11078: waveform_sig_loopback =5506;
11079: waveform_sig_loopback =7313;
11080: waveform_sig_loopback =8010;
11081: waveform_sig_loopback =5768;
11082: waveform_sig_loopback =8709;
11083: waveform_sig_loopback =5226;
11084: waveform_sig_loopback =5347;
11085: waveform_sig_loopback =9685;
11086: waveform_sig_loopback =6967;
11087: waveform_sig_loopback =6227;
11088: waveform_sig_loopback =5703;
11089: waveform_sig_loopback =7892;
11090: waveform_sig_loopback =8480;
11091: waveform_sig_loopback =6041;
11092: waveform_sig_loopback =6497;
11093: waveform_sig_loopback =7696;
11094: waveform_sig_loopback =6732;
11095: waveform_sig_loopback =7854;
11096: waveform_sig_loopback =5883;
11097: waveform_sig_loopback =7594;
11098: waveform_sig_loopback =7826;
11099: waveform_sig_loopback =5992;
11100: waveform_sig_loopback =7755;
11101: waveform_sig_loopback =6871;
11102: waveform_sig_loopback =7287;
11103: waveform_sig_loopback =6566;
11104: waveform_sig_loopback =8069;
11105: waveform_sig_loopback =6780;
11106: waveform_sig_loopback =6539;
11107: waveform_sig_loopback =8007;
11108: waveform_sig_loopback =7170;
11109: waveform_sig_loopback =6531;
11110: waveform_sig_loopback =7358;
11111: waveform_sig_loopback =8265;
11112: waveform_sig_loopback =5770;
11113: waveform_sig_loopback =7397;
11114: waveform_sig_loopback =8617;
11115: waveform_sig_loopback =5909;
11116: waveform_sig_loopback =6765;
11117: waveform_sig_loopback =8326;
11118: waveform_sig_loopback =7386;
11119: waveform_sig_loopback =6076;
11120: waveform_sig_loopback =7322;
11121: waveform_sig_loopback =8765;
11122: waveform_sig_loopback =5786;
11123: waveform_sig_loopback =8927;
11124: waveform_sig_loopback =5643;
11125: waveform_sig_loopback =5354;
11126: waveform_sig_loopback =10345;
11127: waveform_sig_loopback =7009;
11128: waveform_sig_loopback =6105;
11129: waveform_sig_loopback =6536;
11130: waveform_sig_loopback =7797;
11131: waveform_sig_loopback =8595;
11132: waveform_sig_loopback =6307;
11133: waveform_sig_loopback =6506;
11134: waveform_sig_loopback =8006;
11135: waveform_sig_loopback =6813;
11136: waveform_sig_loopback =7835;
11137: waveform_sig_loopback =6217;
11138: waveform_sig_loopback =7703;
11139: waveform_sig_loopback =7706;
11140: waveform_sig_loopback =6319;
11141: waveform_sig_loopback =7757;
11142: waveform_sig_loopback =6967;
11143: waveform_sig_loopback =7456;
11144: waveform_sig_loopback =6420;
11145: waveform_sig_loopback =8170;
11146: waveform_sig_loopback =6881;
11147: waveform_sig_loopback =6249;
11148: waveform_sig_loopback =8267;
11149: waveform_sig_loopback =7002;
11150: waveform_sig_loopback =6273;
11151: waveform_sig_loopback =7854;
11152: waveform_sig_loopback =7623;
11153: waveform_sig_loopback =5876;
11154: waveform_sig_loopback =7489;
11155: waveform_sig_loopback =8063;
11156: waveform_sig_loopback =6239;
11157: waveform_sig_loopback =6484;
11158: waveform_sig_loopback =8162;
11159: waveform_sig_loopback =7457;
11160: waveform_sig_loopback =5513;
11161: waveform_sig_loopback =7495;
11162: waveform_sig_loopback =8496;
11163: waveform_sig_loopback =5285;
11164: waveform_sig_loopback =9254;
11165: waveform_sig_loopback =4934;
11166: waveform_sig_loopback =5358;
11167: waveform_sig_loopback =10346;
11168: waveform_sig_loopback =6305;
11169: waveform_sig_loopback =6094;
11170: waveform_sig_loopback =6230;
11171: waveform_sig_loopback =7505;
11172: waveform_sig_loopback =8502;
11173: waveform_sig_loopback =5785;
11174: waveform_sig_loopback =6283;
11175: waveform_sig_loopback =7724;
11176: waveform_sig_loopback =6440;
11177: waveform_sig_loopback =7370;
11178: waveform_sig_loopback =5986;
11179: waveform_sig_loopback =7313;
11180: waveform_sig_loopback =7267;
11181: waveform_sig_loopback =6101;
11182: waveform_sig_loopback =7033;
11183: waveform_sig_loopback =6788;
11184: waveform_sig_loopback =7030;
11185: waveform_sig_loopback =5708;
11186: waveform_sig_loopback =8198;
11187: waveform_sig_loopback =5929;
11188: waveform_sig_loopback =6093;
11189: waveform_sig_loopback =8005;
11190: waveform_sig_loopback =5936;
11191: waveform_sig_loopback =6328;
11192: waveform_sig_loopback =7104;
11193: waveform_sig_loopback =7021;
11194: waveform_sig_loopback =5692;
11195: waveform_sig_loopback =6620;
11196: waveform_sig_loopback =7717;
11197: waveform_sig_loopback =5561;
11198: waveform_sig_loopback =5767;
11199: waveform_sig_loopback =7930;
11200: waveform_sig_loopback =6538;
11201: waveform_sig_loopback =4914;
11202: waveform_sig_loopback =7176;
11203: waveform_sig_loopback =7479;
11204: waveform_sig_loopback =4812;
11205: waveform_sig_loopback =8616;
11206: waveform_sig_loopback =3986;
11207: waveform_sig_loopback =5028;
11208: waveform_sig_loopback =9551;
11209: waveform_sig_loopback =5466;
11210: waveform_sig_loopback =5448;
11211: waveform_sig_loopback =5458;
11212: waveform_sig_loopback =6701;
11213: waveform_sig_loopback =7930;
11214: waveform_sig_loopback =4796;
11215: waveform_sig_loopback =5524;
11216: waveform_sig_loopback =7126;
11217: waveform_sig_loopback =5332;
11218: waveform_sig_loopback =6883;
11219: waveform_sig_loopback =5046;
11220: waveform_sig_loopback =6290;
11221: waveform_sig_loopback =6745;
11222: waveform_sig_loopback =4955;
11223: waveform_sig_loopback =6217;
11224: waveform_sig_loopback =6165;
11225: waveform_sig_loopback =5599;
11226: waveform_sig_loopback =5337;
11227: waveform_sig_loopback =7118;
11228: waveform_sig_loopback =4744;
11229: waveform_sig_loopback =5651;
11230: waveform_sig_loopback =6495;
11231: waveform_sig_loopback =5350;
11232: waveform_sig_loopback =5272;
11233: waveform_sig_loopback =5954;
11234: waveform_sig_loopback =6261;
11235: waveform_sig_loopback =4344;
11236: waveform_sig_loopback =5806;
11237: waveform_sig_loopback =6661;
11238: waveform_sig_loopback =4468;
11239: waveform_sig_loopback =4722;
11240: waveform_sig_loopback =6724;
11241: waveform_sig_loopback =5565;
11242: waveform_sig_loopback =3760;
11243: waveform_sig_loopback =6324;
11244: waveform_sig_loopback =5860;
11245: waveform_sig_loopback =4082;
11246: waveform_sig_loopback =7744;
11247: waveform_sig_loopback =2166;
11248: waveform_sig_loopback =4467;
11249: waveform_sig_loopback =8188;
11250: waveform_sig_loopback =4343;
11251: waveform_sig_loopback =4431;
11252: waveform_sig_loopback =3892;
11253: waveform_sig_loopback =5954;
11254: waveform_sig_loopback =6636;
11255: waveform_sig_loopback =3161;
11256: waveform_sig_loopback =4825;
11257: waveform_sig_loopback =5599;
11258: waveform_sig_loopback =4175;
11259: waveform_sig_loopback =5741;
11260: waveform_sig_loopback =3349;
11261: waveform_sig_loopback =5565;
11262: waveform_sig_loopback =5257;
11263: waveform_sig_loopback =3440;
11264: waveform_sig_loopback =5302;
11265: waveform_sig_loopback =4564;
11266: waveform_sig_loopback =4361;
11267: waveform_sig_loopback =4119;
11268: waveform_sig_loopback =5461;
11269: waveform_sig_loopback =3675;
11270: waveform_sig_loopback =4195;
11271: waveform_sig_loopback =5024;
11272: waveform_sig_loopback =4092;
11273: waveform_sig_loopback =3805;
11274: waveform_sig_loopback =4678;
11275: waveform_sig_loopback =4792;
11276: waveform_sig_loopback =2915;
11277: waveform_sig_loopback =4506;
11278: waveform_sig_loopback =5285;
11279: waveform_sig_loopback =2780;
11280: waveform_sig_loopback =3552;
11281: waveform_sig_loopback =5579;
11282: waveform_sig_loopback =3576;
11283: waveform_sig_loopback =2586;
11284: waveform_sig_loopback =4935;
11285: waveform_sig_loopback =4362;
11286: waveform_sig_loopback =2812;
11287: waveform_sig_loopback =5719;
11288: waveform_sig_loopback =867;
11289: waveform_sig_loopback =3414;
11290: waveform_sig_loopback =6075;
11291: waveform_sig_loopback =3085;
11292: waveform_sig_loopback =2812;
11293: waveform_sig_loopback =2316;
11294: waveform_sig_loopback =4824;
11295: waveform_sig_loopback =4530;
11296: waveform_sig_loopback =1972;
11297: waveform_sig_loopback =3362;
11298: waveform_sig_loopback =3592;
11299: waveform_sig_loopback =3108;
11300: waveform_sig_loopback =3864;
11301: waveform_sig_loopback =1793;
11302: waveform_sig_loopback =4238;
11303: waveform_sig_loopback =3222;
11304: waveform_sig_loopback =2221;
11305: waveform_sig_loopback =3624;
11306: waveform_sig_loopback =2724;
11307: waveform_sig_loopback =2963;
11308: waveform_sig_loopback =2374;
11309: waveform_sig_loopback =3885;
11310: waveform_sig_loopback =1951;
11311: waveform_sig_loopback =2609;
11312: waveform_sig_loopback =3358;
11313: waveform_sig_loopback =2512;
11314: waveform_sig_loopback =1961;
11315: waveform_sig_loopback =3112;
11316: waveform_sig_loopback =3253;
11317: waveform_sig_loopback =910;
11318: waveform_sig_loopback =3176;
11319: waveform_sig_loopback =3418;
11320: waveform_sig_loopback =909;
11321: waveform_sig_loopback =2252;
11322: waveform_sig_loopback =3460;
11323: waveform_sig_loopback =2003;
11324: waveform_sig_loopback =993;
11325: waveform_sig_loopback =2971;
11326: waveform_sig_loopback =2866;
11327: waveform_sig_loopback =997;
11328: waveform_sig_loopback =3915;
11329: waveform_sig_loopback =-748;
11330: waveform_sig_loopback =1579;
11331: waveform_sig_loopback =4501;
11332: waveform_sig_loopback =1297;
11333: waveform_sig_loopback =722;
11334: waveform_sig_loopback =997;
11335: waveform_sig_loopback =2863;
11336: waveform_sig_loopback =2648;
11337: waveform_sig_loopback =395;
11338: waveform_sig_loopback =1419;
11339: waveform_sig_loopback =1964;
11340: waveform_sig_loopback =1354;
11341: waveform_sig_loopback =1889;
11342: waveform_sig_loopback =236;
11343: waveform_sig_loopback =2361;
11344: waveform_sig_loopback =1255;
11345: waveform_sig_loopback =646;
11346: waveform_sig_loopback =1678;
11347: waveform_sig_loopback =931;
11348: waveform_sig_loopback =1201;
11349: waveform_sig_loopback =521;
11350: waveform_sig_loopback =2123;
11351: waveform_sig_loopback =114;
11352: waveform_sig_loopback =665;
11353: waveform_sig_loopback =1735;
11354: waveform_sig_loopback =551;
11355: waveform_sig_loopback =-52;
11356: waveform_sig_loopback =1714;
11357: waveform_sig_loopback =958;
11358: waveform_sig_loopback =-786;
11359: waveform_sig_loopback =1547;
11360: waveform_sig_loopback =1206;
11361: waveform_sig_loopback =-655;
11362: waveform_sig_loopback =320;
11363: waveform_sig_loopback =1560;
11364: waveform_sig_loopback =297;
11365: waveform_sig_loopback =-1152;
11366: waveform_sig_loopback =1309;
11367: waveform_sig_loopback =965;
11368: waveform_sig_loopback =-1068;
11369: waveform_sig_loopback =2197;
11370: waveform_sig_loopback =-2842;
11371: waveform_sig_loopback =-235;
11372: waveform_sig_loopback =2761;
11373: waveform_sig_loopback =-852;
11374: waveform_sig_loopback =-1160;
11375: waveform_sig_loopback =-642;
11376: waveform_sig_loopback =672;
11377: waveform_sig_loopback =951;
11378: waveform_sig_loopback =-1629;
11379: waveform_sig_loopback =-627;
11380: waveform_sig_loopback =335;
11381: waveform_sig_loopback =-811;
11382: waveform_sig_loopback =-45;
11383: waveform_sig_loopback =-1493;
11384: waveform_sig_loopback =277;
11385: waveform_sig_loopback =-556;
11386: waveform_sig_loopback =-1260;
11387: waveform_sig_loopback =-313;
11388: waveform_sig_loopback =-818;
11389: waveform_sig_loopback =-818;
11390: waveform_sig_loopback =-1345;
11391: waveform_sig_loopback =353;
11392: waveform_sig_loopback =-1932;
11393: waveform_sig_loopback =-1193;
11394: waveform_sig_loopback =74;
11395: waveform_sig_loopback =-1662;
11396: waveform_sig_loopback =-1759;
11397: waveform_sig_loopback =-42;
11398: waveform_sig_loopback =-1376;
11399: waveform_sig_loopback =-2269;
11400: waveform_sig_loopback =-513;
11401: waveform_sig_loopback =-860;
11402: waveform_sig_loopback =-2268;
11403: waveform_sig_loopback =-1920;
11404: waveform_sig_loopback =-24;
11405: waveform_sig_loopback =-1714;
11406: waveform_sig_loopback =-3298;
11407: waveform_sig_loopback =12;
11408: waveform_sig_loopback =-1430;
11409: waveform_sig_loopback =-2768;
11410: waveform_sig_loopback =543;
11411: waveform_sig_loopback =-5208;
11412: waveform_sig_loopback =-1500;
11413: waveform_sig_loopback =674;
11414: waveform_sig_loopback =-2932;
11415: waveform_sig_loopback =-2739;
11416: waveform_sig_loopback =-2700;
11417: waveform_sig_loopback =-1099;
11418: waveform_sig_loopback =-801;
11419: waveform_sig_loopback =-3790;
11420: waveform_sig_loopback =-2231;
11421: waveform_sig_loopback =-1521;
11422: waveform_sig_loopback =-2790;
11423: waveform_sig_loopback =-1733;
11424: waveform_sig_loopback =-3454;
11425: waveform_sig_loopback =-1537;
11426: waveform_sig_loopback =-2349;
11427: waveform_sig_loopback =-3136;
11428: waveform_sig_loopback =-2203;
11429: waveform_sig_loopback =-2501;
11430: waveform_sig_loopback =-2850;
11431: waveform_sig_loopback =-3064;
11432: waveform_sig_loopback =-1376;
11433: waveform_sig_loopback =-4143;
11434: waveform_sig_loopback =-2593;
11435: waveform_sig_loopback =-1916;
11436: waveform_sig_loopback =-3716;
11437: waveform_sig_loopback =-3090;
11438: waveform_sig_loopback =-2245;
11439: waveform_sig_loopback =-3079;
11440: waveform_sig_loopback =-3924;
11441: waveform_sig_loopback =-2628;
11442: waveform_sig_loopback =-2217;
11443: waveform_sig_loopback =-4423;
11444: waveform_sig_loopback =-3651;
11445: waveform_sig_loopback =-1461;
11446: waveform_sig_loopback =-4029;
11447: waveform_sig_loopback =-4723;
11448: waveform_sig_loopback =-1707;
11449: waveform_sig_loopback =-3609;
11450: waveform_sig_loopback =-3999;
11451: waveform_sig_loopback =-1586;
11452: waveform_sig_loopback =-7093;
11453: waveform_sig_loopback =-2753;
11454: waveform_sig_loopback =-1461;
11455: waveform_sig_loopback =-4527;
11456: waveform_sig_loopback =-4451;
11457: waveform_sig_loopback =-4588;
11458: waveform_sig_loopback =-2485;
11459: waveform_sig_loopback =-2662;
11460: waveform_sig_loopback =-5678;
11461: waveform_sig_loopback =-3634;
11462: waveform_sig_loopback =-3455;
11463: waveform_sig_loopback =-4418;
11464: waveform_sig_loopback =-3314;
11465: waveform_sig_loopback =-5365;
11466: waveform_sig_loopback =-3014;
11467: waveform_sig_loopback =-4000;
11468: waveform_sig_loopback =-5015;
11469: waveform_sig_loopback =-3700;
11470: waveform_sig_loopback =-4130;
11471: waveform_sig_loopback =-4789;
11472: waveform_sig_loopback =-4279;
11473: waveform_sig_loopback =-3356;
11474: waveform_sig_loopback =-5813;
11475: waveform_sig_loopback =-3800;
11476: waveform_sig_loopback =-4112;
11477: waveform_sig_loopback =-4886;
11478: waveform_sig_loopback =-4871;
11479: waveform_sig_loopback =-4052;
11480: waveform_sig_loopback =-4191;
11481: waveform_sig_loopback =-6076;
11482: waveform_sig_loopback =-3812;
11483: waveform_sig_loopback =-3816;
11484: waveform_sig_loopback =-6391;
11485: waveform_sig_loopback =-4673;
11486: waveform_sig_loopback =-3376;
11487: waveform_sig_loopback =-5565;
11488: waveform_sig_loopback =-6042;
11489: waveform_sig_loopback =-3439;
11490: waveform_sig_loopback =-5039;
11491: waveform_sig_loopback =-5458;
11492: waveform_sig_loopback =-3225;
11493: waveform_sig_loopback =-8631;
11494: waveform_sig_loopback =-3988;
11495: waveform_sig_loopback =-3098;
11496: waveform_sig_loopback =-6127;
11497: waveform_sig_loopback =-5832;
11498: waveform_sig_loopback =-6162;
11499: waveform_sig_loopback =-3672;
11500: waveform_sig_loopback =-4386;
11501: waveform_sig_loopback =-7233;
11502: waveform_sig_loopback =-4581;
11503: waveform_sig_loopback =-5405;
11504: waveform_sig_loopback =-5481;
11505: waveform_sig_loopback =-4811;
11506: waveform_sig_loopback =-7016;
11507: waveform_sig_loopback =-3899;
11508: waveform_sig_loopback =-5901;
11509: waveform_sig_loopback =-6205;
11510: waveform_sig_loopback =-4798;
11511: waveform_sig_loopback =-5959;
11512: waveform_sig_loopback =-5762;
11513: waveform_sig_loopback =-5741;
11514: waveform_sig_loopback =-4947;
11515: waveform_sig_loopback =-6693;
11516: waveform_sig_loopback =-5588;
11517: waveform_sig_loopback =-5245;
11518: waveform_sig_loopback =-6150;
11519: waveform_sig_loopback =-6451;
11520: waveform_sig_loopback =-4916;
11521: waveform_sig_loopback =-5866;
11522: waveform_sig_loopback =-7297;
11523: waveform_sig_loopback =-4836;
11524: waveform_sig_loopback =-5383;
11525: waveform_sig_loopback =-7593;
11526: waveform_sig_loopback =-5777;
11527: waveform_sig_loopback =-4704;
11528: waveform_sig_loopback =-6879;
11529: waveform_sig_loopback =-7127;
11530: waveform_sig_loopback =-4739;
11531: waveform_sig_loopback =-6256;
11532: waveform_sig_loopback =-6466;
11533: waveform_sig_loopback =-4688;
11534: waveform_sig_loopback =-9657;
11535: waveform_sig_loopback =-5075;
11536: waveform_sig_loopback =-4495;
11537: waveform_sig_loopback =-6880;
11538: waveform_sig_loopback =-7365;
11539: waveform_sig_loopback =-7011;
11540: waveform_sig_loopback =-4647;
11541: waveform_sig_loopback =-5930;
11542: waveform_sig_loopback =-7820;
11543: waveform_sig_loopback =-5959;
11544: waveform_sig_loopback =-6516;
11545: waveform_sig_loopback =-6102;
11546: waveform_sig_loopback =-6418;
11547: waveform_sig_loopback =-7577;
11548: waveform_sig_loopback =-5002;
11549: waveform_sig_loopback =-7303;
11550: waveform_sig_loopback =-6646;
11551: waveform_sig_loopback =-6285;
11552: waveform_sig_loopback =-6731;
11553: waveform_sig_loopback =-6604;
11554: waveform_sig_loopback =-7004;
11555: waveform_sig_loopback =-5579;
11556: waveform_sig_loopback =-7885;
11557: waveform_sig_loopback =-6415;
11558: waveform_sig_loopback =-6048;
11559: waveform_sig_loopback =-7260;
11560: waveform_sig_loopback =-7172;
11561: waveform_sig_loopback =-5750;
11562: waveform_sig_loopback =-6839;
11563: waveform_sig_loopback =-8084;
11564: waveform_sig_loopback =-5549;
11565: waveform_sig_loopback =-6467;
11566: waveform_sig_loopback =-8340;
11567: waveform_sig_loopback =-6315;
11568: waveform_sig_loopback =-5852;
11569: waveform_sig_loopback =-7453;
11570: waveform_sig_loopback =-7953;
11571: waveform_sig_loopback =-5539;
11572: waveform_sig_loopback =-6832;
11573: waveform_sig_loopback =-7473;
11574: waveform_sig_loopback =-5373;
11575: waveform_sig_loopback =-10216;
11576: waveform_sig_loopback =-5986;
11577: waveform_sig_loopback =-4848;
11578: waveform_sig_loopback =-8009;
11579: waveform_sig_loopback =-8020;
11580: waveform_sig_loopback =-7222;
11581: waveform_sig_loopback =-5850;
11582: waveform_sig_loopback =-6262;
11583: waveform_sig_loopback =-8532;
11584: waveform_sig_loopback =-6773;
11585: waveform_sig_loopback =-6761;
11586: waveform_sig_loopback =-7091;
11587: waveform_sig_loopback =-6913;
11588: waveform_sig_loopback =-8108;
11589: waveform_sig_loopback =-5922;
11590: waveform_sig_loopback =-7449;
11591: waveform_sig_loopback =-7346;
11592: waveform_sig_loopback =-7102;
11593: waveform_sig_loopback =-7108;
11594: waveform_sig_loopback =-7184;
11595: waveform_sig_loopback =-7316;
11596: waveform_sig_loopback =-6249;
11597: waveform_sig_loopback =-8478;
11598: waveform_sig_loopback =-6667;
11599: waveform_sig_loopback =-6453;
11600: waveform_sig_loopback =-8019;
11601: waveform_sig_loopback =-7546;
11602: waveform_sig_loopback =-5953;
11603: waveform_sig_loopback =-7735;
11604: waveform_sig_loopback =-8165;
11605: waveform_sig_loopback =-6018;
11606: waveform_sig_loopback =-7023;
11607: waveform_sig_loopback =-8376;
11608: waveform_sig_loopback =-7154;
11609: waveform_sig_loopback =-5881;
11610: waveform_sig_loopback =-7767;
11611: waveform_sig_loopback =-8713;
11612: waveform_sig_loopback =-5365;
11613: waveform_sig_loopback =-7625;
11614: waveform_sig_loopback =-7429;
11615: waveform_sig_loopback =-5572;
11616: waveform_sig_loopback =-11254;
11617: waveform_sig_loopback =-5483;
11618: waveform_sig_loopback =-5296;
11619: waveform_sig_loopback =-8483;
11620: waveform_sig_loopback =-7885;
11621: waveform_sig_loopback =-7868;
11622: waveform_sig_loopback =-5882;
11623: waveform_sig_loopback =-6443;
11624: waveform_sig_loopback =-8988;
11625: waveform_sig_loopback =-6646;
11626: waveform_sig_loopback =-7144;
11627: waveform_sig_loopback =-7327;
11628: waveform_sig_loopback =-6935;
11629: waveform_sig_loopback =-8134;
11630: waveform_sig_loopback =-6088;
11631: waveform_sig_loopback =-7622;
11632: waveform_sig_loopback =-7604;
11633: waveform_sig_loopback =-6954;
11634: waveform_sig_loopback =-6856;
11635: waveform_sig_loopback =-7852;
11636: waveform_sig_loopback =-7177;
11637: waveform_sig_loopback =-6082;
11638: waveform_sig_loopback =-8705;
11639: waveform_sig_loopback =-6463;
11640: waveform_sig_loopback =-6799;
11641: waveform_sig_loopback =-7855;
11642: waveform_sig_loopback =-7114;
11643: waveform_sig_loopback =-6504;
11644: waveform_sig_loopback =-7376;
11645: waveform_sig_loopback =-7954;
11646: waveform_sig_loopback =-6243;
11647: waveform_sig_loopback =-6642;
11648: waveform_sig_loopback =-8547;
11649: waveform_sig_loopback =-6742;
11650: waveform_sig_loopback =-5685;
11651: waveform_sig_loopback =-8155;
11652: waveform_sig_loopback =-8047;
11653: waveform_sig_loopback =-5118;
11654: waveform_sig_loopback =-7826;
11655: waveform_sig_loopback =-6819;
11656: waveform_sig_loopback =-5733;
11657: waveform_sig_loopback =-10884;
11658: waveform_sig_loopback =-4817;
11659: waveform_sig_loopback =-5657;
11660: waveform_sig_loopback =-8081;
11661: waveform_sig_loopback =-7559;
11662: waveform_sig_loopback =-7680;
11663: waveform_sig_loopback =-5210;
11664: waveform_sig_loopback =-6458;
11665: waveform_sig_loopback =-8732;
11666: waveform_sig_loopback =-5937;
11667: waveform_sig_loopback =-7102;
11668: waveform_sig_loopback =-6713;
11669: waveform_sig_loopback =-6618;
11670: waveform_sig_loopback =-7971;
11671: waveform_sig_loopback =-5365;
11672: waveform_sig_loopback =-7328;
11673: waveform_sig_loopback =-7186;
11674: waveform_sig_loopback =-6393;
11675: waveform_sig_loopback =-6602;
11676: waveform_sig_loopback =-7385;
11677: waveform_sig_loopback =-6307;
11678: waveform_sig_loopback =-6077;
11679: waveform_sig_loopback =-8038;
11680: waveform_sig_loopback =-5799;
11681: waveform_sig_loopback =-6649;
11682: waveform_sig_loopback =-6911;
11683: waveform_sig_loopback =-6946;
11684: waveform_sig_loopback =-5791;
11685: waveform_sig_loopback =-6598;
11686: waveform_sig_loopback =-7779;
11687: waveform_sig_loopback =-5240;
11688: waveform_sig_loopback =-6265;
11689: waveform_sig_loopback =-8019;
11690: waveform_sig_loopback =-5857;
11691: waveform_sig_loopback =-5357;
11692: waveform_sig_loopback =-7451;
11693: waveform_sig_loopback =-7244;
11694: waveform_sig_loopback =-4636;
11695: waveform_sig_loopback =-7233;
11696: waveform_sig_loopback =-5923;
11697: waveform_sig_loopback =-5452;
11698: waveform_sig_loopback =-10029;
11699: waveform_sig_loopback =-3915;
11700: waveform_sig_loopback =-5203;
11701: waveform_sig_loopback =-7122;
11702: waveform_sig_loopback =-7038;
11703: waveform_sig_loopback =-6782;
11704: waveform_sig_loopback =-4203;
11705: waveform_sig_loopback =-6093;
11706: waveform_sig_loopback =-7736;
11707: waveform_sig_loopback =-5049;
11708: waveform_sig_loopback =-6564;
11709: waveform_sig_loopback =-5532;
11710: waveform_sig_loopback =-6126;
11711: waveform_sig_loopback =-7068;
11712: waveform_sig_loopback =-4300;
11713: waveform_sig_loopback =-6898;
11714: waveform_sig_loopback =-5987;
11715: waveform_sig_loopback =-5521;
11716: waveform_sig_loopback =-5938;
11717: waveform_sig_loopback =-6202;
11718: waveform_sig_loopback =-5583;
11719: waveform_sig_loopback =-5167;
11720: waveform_sig_loopback =-6895;
11721: waveform_sig_loopback =-5117;
11722: waveform_sig_loopback =-5440;
11723: waveform_sig_loopback =-6078;
11724: waveform_sig_loopback =-6019;
11725: waveform_sig_loopback =-4618;
11726: waveform_sig_loopback =-5894;
11727: waveform_sig_loopback =-6664;
11728: waveform_sig_loopback =-4100;
11729: waveform_sig_loopback =-5420;
11730: waveform_sig_loopback =-6954;
11731: waveform_sig_loopback =-4647;
11732: waveform_sig_loopback =-4434;
11733: waveform_sig_loopback =-6386;
11734: waveform_sig_loopback =-5949;
11735: waveform_sig_loopback =-3750;
11736: waveform_sig_loopback =-6040;
11737: waveform_sig_loopback =-4685;
11738: waveform_sig_loopback =-4620;
11739: waveform_sig_loopback =-8488;
11740: waveform_sig_loopback =-2996;
11741: waveform_sig_loopback =-4008;
11742: waveform_sig_loopback =-5801;
11743: waveform_sig_loopback =-6231;
11744: waveform_sig_loopback =-5142;
11745: waveform_sig_loopback =-3272;
11746: waveform_sig_loopback =-4944;
11747: waveform_sig_loopback =-6254;
11748: waveform_sig_loopback =-4194;
11749: waveform_sig_loopback =-5088;
11750: waveform_sig_loopback =-4314;
11751: waveform_sig_loopback =-5098;
11752: waveform_sig_loopback =-5445;
11753: waveform_sig_loopback =-3235;
11754: waveform_sig_loopback =-5663;
11755: waveform_sig_loopback =-4479;
11756: waveform_sig_loopback =-4431;
11757: waveform_sig_loopback =-4542;
11758: waveform_sig_loopback =-4881;
11759: waveform_sig_loopback =-4318;
11760: waveform_sig_loopback =-3802;
11761: waveform_sig_loopback =-5556;
11762: waveform_sig_loopback =-3819;
11763: waveform_sig_loopback =-3938;
11764: waveform_sig_loopback =-4864;
11765: waveform_sig_loopback =-4606;
11766: waveform_sig_loopback =-2990;
11767: waveform_sig_loopback =-4914;
11768: waveform_sig_loopback =-4973;
11769: waveform_sig_loopback =-2692;
11770: waveform_sig_loopback =-4332;
11771: waveform_sig_loopback =-5225;
11772: waveform_sig_loopback =-3341;
11773: waveform_sig_loopback =-3023;
11774: waveform_sig_loopback =-4872;
11775: waveform_sig_loopback =-4627;
11776: waveform_sig_loopback =-2096;
11777: waveform_sig_loopback =-4675;
11778: waveform_sig_loopback =-3214;
11779: waveform_sig_loopback =-3166;
11780: waveform_sig_loopback =-7022;
11781: waveform_sig_loopback =-1396;
11782: waveform_sig_loopback =-2409;
11783: waveform_sig_loopback =-4591;
11784: waveform_sig_loopback =-4619;
11785: waveform_sig_loopback =-3364;
11786: waveform_sig_loopback =-2012;
11787: waveform_sig_loopback =-3244;
11788: waveform_sig_loopback =-4824;
11789: waveform_sig_loopback =-2613;
11790: waveform_sig_loopback =-3307;
11791: waveform_sig_loopback =-3012;
11792: waveform_sig_loopback =-3412;
11793: waveform_sig_loopback =-3733;
11794: waveform_sig_loopback =-1886;
11795: waveform_sig_loopback =-3911;
11796: waveform_sig_loopback =-2959;
11797: waveform_sig_loopback =-2855;
11798: waveform_sig_loopback =-2810;
11799: waveform_sig_loopback =-3417;
11800: waveform_sig_loopback =-2549;
11801: waveform_sig_loopback =-2167;
11802: waveform_sig_loopback =-4042;
11803: waveform_sig_loopback =-2076;
11804: waveform_sig_loopback =-2179;
11805: waveform_sig_loopback =-3483;
11806: waveform_sig_loopback =-2637;
11807: waveform_sig_loopback =-1433;
11808: waveform_sig_loopback =-3426;
11809: waveform_sig_loopback =-2888;
11810: waveform_sig_loopback =-1317;
11811: waveform_sig_loopback =-2507;
11812: waveform_sig_loopback =-3432;
11813: waveform_sig_loopback =-1808;
11814: waveform_sig_loopback =-1083;
11815: waveform_sig_loopback =-3421;
11816: waveform_sig_loopback =-2813;
11817: waveform_sig_loopback =-156;
11818: waveform_sig_loopback =-3291;
11819: waveform_sig_loopback =-1186;
11820: waveform_sig_loopback =-1608;
11821: waveform_sig_loopback =-5370;
11822: waveform_sig_loopback =727;
11823: waveform_sig_loopback =-942;
11824: waveform_sig_loopback =-2919;
11825: waveform_sig_loopback =-2567;
11826: waveform_sig_loopback =-1779;
11827: waveform_sig_loopback =-116;
11828: waveform_sig_loopback =-1435;
11829: waveform_sig_loopback =-3218;
11830: waveform_sig_loopback =-613;
11831: waveform_sig_loopback =-1630;
11832: waveform_sig_loopback =-1255;
11833: waveform_sig_loopback =-1503;
11834: waveform_sig_loopback =-1981;
11835: waveform_sig_loopback =-13;
11836: waveform_sig_loopback =-1985;
11837: waveform_sig_loopback =-1304;
11838: waveform_sig_loopback =-928;
11839: waveform_sig_loopback =-917;
11840: waveform_sig_loopback =-1797;
11841: waveform_sig_loopback =-428;
11842: waveform_sig_loopback =-523;
11843: waveform_sig_loopback =-2250;
11844: waveform_sig_loopback =48;
11845: waveform_sig_loopback =-671;
11846: waveform_sig_loopback =-1521;
11847: waveform_sig_loopback =-643;
11848: waveform_sig_loopback =143;
11849: waveform_sig_loopback =-1370;
11850: waveform_sig_loopback =-1111;
11851: waveform_sig_loopback =545;
11852: waveform_sig_loopback =-557;
11853: waveform_sig_loopback =-1779;
11854: waveform_sig_loopback =275;
11855: waveform_sig_loopback =796;
11856: waveform_sig_loopback =-1758;
11857: waveform_sig_loopback =-729;
11858: waveform_sig_loopback =1698;
11859: waveform_sig_loopback =-1633;
11860: waveform_sig_loopback =1078;
11861: waveform_sig_loopback =-96;
11862: waveform_sig_loopback =-3425;
11863: waveform_sig_loopback =2982;
11864: waveform_sig_loopback =486;
11865: waveform_sig_loopback =-842;
11866: waveform_sig_loopback =-633;
11867: waveform_sig_loopback =-108;
11868: waveform_sig_loopback =2099;
11869: waveform_sig_loopback =25;
11870: waveform_sig_loopback =-1260;
11871: waveform_sig_loopback =1545;
11872: waveform_sig_loopback =-167;
11873: waveform_sig_loopback =941;
11874: waveform_sig_loopback =190;
11875: waveform_sig_loopback =-182;
11876: waveform_sig_loopback =2093;
11877: waveform_sig_loopback =-396;
11878: waveform_sig_loopback =737;
11879: waveform_sig_loopback =918;
11880: waveform_sig_loopback =843;
11881: waveform_sig_loopback =167;
11882: waveform_sig_loopback =1539;
11883: waveform_sig_loopback =1141;
11884: waveform_sig_loopback =-292;
11885: waveform_sig_loopback =2076;
11886: waveform_sig_loopback =1019;
11887: waveform_sig_loopback =551;
11888: waveform_sig_loopback =1212;
11889: waveform_sig_loopback =1882;
11890: waveform_sig_loopback =798;
11891: waveform_sig_loopback =589;
11892: waveform_sig_loopback =2591;
11893: waveform_sig_loopback =1336;
11894: waveform_sig_loopback =-84;
11895: waveform_sig_loopback =2640;
11896: waveform_sig_loopback =2362;
11897: waveform_sig_loopback =32;
11898: waveform_sig_loopback =1633;
11899: waveform_sig_loopback =3143;
11900: waveform_sig_loopback =396;
11901: waveform_sig_loopback =3192;
11902: waveform_sig_loopback =1273;
11903: waveform_sig_loopback =-1048;
11904: waveform_sig_loopback =4726;
11905: waveform_sig_loopback =2295;
11906: waveform_sig_loopback =1247;
11907: waveform_sig_loopback =868;
11908: waveform_sig_loopback =2097;
11909: waveform_sig_loopback =4033;
11910: waveform_sig_loopback =1609;
11911: waveform_sig_loopback =887;
11912: waveform_sig_loopback =3300;
11913: waveform_sig_loopback =1697;
11914: waveform_sig_loopback =3094;
11915: waveform_sig_loopback =1775;
11916: waveform_sig_loopback =1926;
11917: waveform_sig_loopback =3971;
11918: waveform_sig_loopback =1332;
11919: waveform_sig_loopback =2754;
11920: waveform_sig_loopback =2762;
11921: waveform_sig_loopback =2625;
11922: waveform_sig_loopback =2099;
11923: waveform_sig_loopback =3479;
11924: waveform_sig_loopback =2708;
11925: waveform_sig_loopback =1914;
11926: waveform_sig_loopback =3711;
11927: waveform_sig_loopback =2792;
11928: waveform_sig_loopback =2589;
11929: waveform_sig_loopback =2698;
11930: waveform_sig_loopback =4109;
11931: waveform_sig_loopback =2270;
11932: waveform_sig_loopback =2336;
11933: waveform_sig_loopback =4738;
11934: waveform_sig_loopback =2590;
11935: waveform_sig_loopback =1993;
11936: waveform_sig_loopback =4426;
11937: waveform_sig_loopback =3841;
11938: waveform_sig_loopback =1912;
11939: waveform_sig_loopback =3303;
11940: waveform_sig_loopback =4988;
11941: waveform_sig_loopback =2256;
11942: waveform_sig_loopback =4646;
11943: waveform_sig_loopback =2874;
11944: waveform_sig_loopback =1083;
11945: waveform_sig_loopback =6376;
11946: waveform_sig_loopback =3966;
11947: waveform_sig_loopback =2756;
11948: waveform_sig_loopback =2769;
11949: waveform_sig_loopback =3964;
11950: waveform_sig_loopback =5485;
11951: waveform_sig_loopback =3257;
11952: waveform_sig_loopback =2737;
11953: waveform_sig_loopback =5002;
11954: waveform_sig_loopback =3213;
11955: waveform_sig_loopback =4897;
11956: waveform_sig_loopback =3243;
11957: waveform_sig_loopback =3825;
11958: waveform_sig_loopback =5494;
11959: waveform_sig_loopback =2760;
11960: waveform_sig_loopback =4754;
11961: waveform_sig_loopback =4221;
11962: waveform_sig_loopback =4129;
11963: waveform_sig_loopback =3954;
11964: waveform_sig_loopback =4852;
11965: waveform_sig_loopback =4474;
11966: waveform_sig_loopback =3533;
11967: waveform_sig_loopback =5006;
11968: waveform_sig_loopback =4888;
11969: waveform_sig_loopback =3683;
11970: waveform_sig_loopback =4496;
11971: waveform_sig_loopback =5821;
11972: waveform_sig_loopback =3375;
11973: waveform_sig_loopback =4467;
11974: waveform_sig_loopback =5986;
11975: waveform_sig_loopback =4112;
11976: waveform_sig_loopback =3755;
11977: waveform_sig_loopback =5790;
11978: waveform_sig_loopback =5486;
11979: waveform_sig_loopback =3519;
11980: waveform_sig_loopback =4901;
11981: waveform_sig_loopback =6424;
11982: waveform_sig_loopback =3670;
11983: waveform_sig_loopback =6483;
11984: waveform_sig_loopback =4143;
11985: waveform_sig_loopback =2553;
11986: waveform_sig_loopback =7906;
11987: waveform_sig_loopback =5421;
11988: waveform_sig_loopback =4298;
11989: waveform_sig_loopback =3977;
11990: waveform_sig_loopback =5766;
11991: waveform_sig_loopback =6802;
11992: waveform_sig_loopback =4549;
11993: waveform_sig_loopback =4502;
11994: waveform_sig_loopback =5997;
11995: waveform_sig_loopback =5105;
11996: waveform_sig_loopback =6093;
11997: waveform_sig_loopback =4420;
11998: waveform_sig_loopback =5750;
11999: waveform_sig_loopback =6346;
12000: waveform_sig_loopback =4492;
12001: waveform_sig_loopback =6121;
12002: waveform_sig_loopback =5266;
12003: waveform_sig_loopback =6059;
12004: waveform_sig_loopback =4836;
12005: waveform_sig_loopback =6407;
12006: waveform_sig_loopback =5892;
12007: waveform_sig_loopback =4567;
12008: waveform_sig_loopback =6791;
12009: waveform_sig_loopback =5775;
12010: waveform_sig_loopback =5122;
12011: waveform_sig_loopback =6066;
12012: waveform_sig_loopback =6759;
12013: waveform_sig_loopback =4792;
12014: waveform_sig_loopback =5744;
12015: waveform_sig_loopback =7310;
12016: waveform_sig_loopback =5150;
12017: waveform_sig_loopback =5134;
12018: waveform_sig_loopback =7093;
12019: waveform_sig_loopback =6465;
12020: waveform_sig_loopback =4893;
12021: waveform_sig_loopback =5895;
12022: waveform_sig_loopback =7817;
12023: waveform_sig_loopback =4764;
12024: waveform_sig_loopback =7588;
12025: waveform_sig_loopback =5416;
12026: waveform_sig_loopback =3582;
12027: waveform_sig_loopback =9272;
12028: waveform_sig_loopback =6522;
12029: waveform_sig_loopback =5045;
12030: waveform_sig_loopback =5550;
12031: waveform_sig_loopback =6708;
12032: waveform_sig_loopback =7790;
12033: waveform_sig_loopback =5913;
12034: waveform_sig_loopback =5213;
12035: waveform_sig_loopback =7343;
12036: waveform_sig_loopback =6156;
12037: waveform_sig_loopback =6876;
12038: waveform_sig_loopback =5832;
12039: waveform_sig_loopback =6600;
12040: waveform_sig_loopback =7289;
12041: waveform_sig_loopback =5778;
12042: waveform_sig_loopback =6744;
12043: waveform_sig_loopback =6504;
12044: waveform_sig_loopback =6962;
12045: waveform_sig_loopback =5652;
12046: waveform_sig_loopback =7737;
12047: waveform_sig_loopback =6455;
12048: waveform_sig_loopback =5663;
12049: waveform_sig_loopback =7804;
12050: waveform_sig_loopback =6520;
12051: waveform_sig_loopback =6096;
12052: waveform_sig_loopback =6987;
12053: waveform_sig_loopback =7605;
12054: waveform_sig_loopback =5603;
12055: waveform_sig_loopback =6795;
12056: waveform_sig_loopback =7957;
12057: waveform_sig_loopback =6029;
12058: waveform_sig_loopback =6119;
12059: waveform_sig_loopback =7732;
12060: waveform_sig_loopback =7560;
12061: waveform_sig_loopback =5407;
12062: waveform_sig_loopback =6840;
12063: waveform_sig_loopback =8827;
12064: waveform_sig_loopback =5023;
12065: waveform_sig_loopback =8903;
12066: waveform_sig_loopback =5777;
12067: waveform_sig_loopback =4317;
12068: waveform_sig_loopback =10531;
12069: waveform_sig_loopback =6569;
12070: waveform_sig_loopback =6037;
12071: waveform_sig_loopback =6432;
12072: waveform_sig_loopback =7044;
12073: waveform_sig_loopback =8916;
12074: waveform_sig_loopback =6174;
12075: waveform_sig_loopback =6005;
12076: waveform_sig_loopback =8257;
12077: waveform_sig_loopback =6328;
12078: waveform_sig_loopback =7753;
12079: waveform_sig_loopback =6389;
12080: waveform_sig_loopback =7045;
12081: waveform_sig_loopback =8048;
12082: waveform_sig_loopback =6147;
12083: waveform_sig_loopback =7401;
12084: waveform_sig_loopback =7198;
12085: waveform_sig_loopback =7306;
12086: waveform_sig_loopback =6250;
12087: waveform_sig_loopback =8306;
12088: waveform_sig_loopback =6839;
12089: waveform_sig_loopback =6181;
12090: waveform_sig_loopback =8413;
12091: waveform_sig_loopback =6761;
12092: waveform_sig_loopback =6693;
12093: waveform_sig_loopback =7557;
12094: waveform_sig_loopback =7677;
12095: waveform_sig_loopback =6408;
12096: waveform_sig_loopback =6988;
12097: waveform_sig_loopback =8401;
12098: waveform_sig_loopback =6616;
12099: waveform_sig_loopback =6093;
12100: waveform_sig_loopback =8540;
12101: waveform_sig_loopback =7661;
12102: waveform_sig_loopback =5527;
12103: waveform_sig_loopback =7749;
12104: waveform_sig_loopback =8581;
12105: waveform_sig_loopback =5534;
12106: waveform_sig_loopback =9415;
12107: waveform_sig_loopback =5395;
12108: waveform_sig_loopback =5297;
12109: waveform_sig_loopback =10508;
12110: waveform_sig_loopback =6671;
12111: waveform_sig_loopback =6643;
12112: waveform_sig_loopback =6199;
12113: waveform_sig_loopback =7598;
12114: waveform_sig_loopback =9092;
12115: waveform_sig_loopback =6064;
12116: waveform_sig_loopback =6479;
12117: waveform_sig_loopback =8245;
12118: waveform_sig_loopback =6502;
12119: waveform_sig_loopback =8079;
12120: waveform_sig_loopback =6252;
12121: waveform_sig_loopback =7279;
12122: waveform_sig_loopback =8265;
12123: waveform_sig_loopback =6039;
12124: waveform_sig_loopback =7549;
12125: waveform_sig_loopback =7345;
12126: waveform_sig_loopback =7120;
12127: waveform_sig_loopback =6489;
12128: waveform_sig_loopback =8328;
12129: waveform_sig_loopback =6531;
12130: waveform_sig_loopback =6657;
12131: waveform_sig_loopback =8048;
12132: waveform_sig_loopback =6758;
12133: waveform_sig_loopback =6843;
12134: waveform_sig_loopback =7197;
12135: waveform_sig_loopback =7943;
12136: waveform_sig_loopback =6087;
12137: waveform_sig_loopback =6906;
12138: waveform_sig_loopback =8543;
12139: waveform_sig_loopback =6129;
12140: waveform_sig_loopback =6146;
12141: waveform_sig_loopback =8551;
12142: waveform_sig_loopback =7212;
12143: waveform_sig_loopback =5544;
12144: waveform_sig_loopback =7664;
12145: waveform_sig_loopback =8128;
12146: waveform_sig_loopback =5672;
12147: waveform_sig_loopback =9085;
12148: waveform_sig_loopback =4923;
12149: waveform_sig_loopback =5563;
12150: waveform_sig_loopback =9951;
12151: waveform_sig_loopback =6527;
12152: waveform_sig_loopback =6359;
12153: waveform_sig_loopback =5734;
12154: waveform_sig_loopback =7683;
12155: waveform_sig_loopback =8567;
12156: waveform_sig_loopback =5661;
12157: waveform_sig_loopback =6430;
12158: waveform_sig_loopback =7666;
12159: waveform_sig_loopback =6302;
12160: waveform_sig_loopback =7782;
12161: waveform_sig_loopback =5582;
12162: waveform_sig_loopback =7265;
12163: waveform_sig_loopback =7730;
12164: waveform_sig_loopback =5544;
12165: waveform_sig_loopback =7376;
12166: waveform_sig_loopback =6715;
12167: waveform_sig_loopback =6679;
12168: waveform_sig_loopback =6274;
12169: waveform_sig_loopback =7647;
12170: waveform_sig_loopback =6186;
12171: waveform_sig_loopback =6228;
12172: waveform_sig_loopback =7369;
12173: waveform_sig_loopback =6609;
12174: waveform_sig_loopback =6015;
12175: waveform_sig_loopback =6828;
12176: waveform_sig_loopback =7559;
12177: waveform_sig_loopback =5159;
12178: waveform_sig_loopback =6733;
12179: waveform_sig_loopback =7921;
12180: waveform_sig_loopback =5296;
12181: waveform_sig_loopback =5913;
12182: waveform_sig_loopback =7775;
12183: waveform_sig_loopback =6518;
12184: waveform_sig_loopback =5113;
12185: waveform_sig_loopback =6902;
12186: waveform_sig_loopback =7504;
12187: waveform_sig_loopback =5058;
12188: waveform_sig_loopback =8278;
12189: waveform_sig_loopback =4262;
12190: waveform_sig_loopback =4983;
12191: waveform_sig_loopback =9125;
12192: waveform_sig_loopback =5999;
12193: waveform_sig_loopback =5350;
12194: waveform_sig_loopback =5080;
12195: waveform_sig_loopback =7205;
12196: waveform_sig_loopback =7414;
12197: waveform_sig_loopback =5010;
12198: waveform_sig_loopback =5679;
12199: waveform_sig_loopback =6669;
12200: waveform_sig_loopback =5823;
12201: waveform_sig_loopback =6629;
12202: waveform_sig_loopback =4859;
12203: waveform_sig_loopback =6702;
12204: waveform_sig_loopback =6426;
12205: waveform_sig_loopback =4943;
12206: waveform_sig_loopback =6502;
12207: waveform_sig_loopback =5667;
12208: waveform_sig_loopback =5987;
12209: waveform_sig_loopback =5227;
12210: waveform_sig_loopback =6771;
12211: waveform_sig_loopback =5291;
12212: waveform_sig_loopback =5151;
12213: waveform_sig_loopback =6565;
12214: waveform_sig_loopback =5631;
12215: waveform_sig_loopback =4813;
12216: waveform_sig_loopback =6149;
12217: waveform_sig_loopback =6377;
12218: waveform_sig_loopback =4050;
12219: waveform_sig_loopback =6036;
12220: waveform_sig_loopback =6573;
12221: waveform_sig_loopback =4325;
12222: waveform_sig_loopback =5097;
12223: waveform_sig_loopback =6474;
12224: waveform_sig_loopback =5586;
12225: waveform_sig_loopback =3956;
12226: waveform_sig_loopback =5831;
12227: waveform_sig_loopback =6555;
12228: waveform_sig_loopback =3724;
12229: waveform_sig_loopback =7295;
12230: waveform_sig_loopback =3038;
12231: waveform_sig_loopback =3840;
12232: waveform_sig_loopback =8255;
12233: waveform_sig_loopback =4581;
12234: waveform_sig_loopback =4044;
12235: waveform_sig_loopback =4291;
12236: waveform_sig_loopback =5836;
12237: waveform_sig_loopback =6277;
12238: waveform_sig_loopback =3896;
12239: waveform_sig_loopback =4320;
12240: waveform_sig_loopback =5665;
12241: waveform_sig_loopback =4495;
12242: waveform_sig_loopback =5339;
12243: waveform_sig_loopback =3806;
12244: waveform_sig_loopback =5355;
12245: waveform_sig_loopback =5120;
12246: waveform_sig_loopback =3872;
12247: waveform_sig_loopback =5074;
12248: waveform_sig_loopback =4440;
12249: waveform_sig_loopback =4788;
12250: waveform_sig_loopback =3704;
12251: waveform_sig_loopback =5670;
12252: waveform_sig_loopback =3921;
12253: waveform_sig_loopback =3660;
12254: waveform_sig_loopback =5567;
12255: waveform_sig_loopback =3955;
12256: waveform_sig_loopback =3586;
12257: waveform_sig_loopback =5076;
12258: waveform_sig_loopback =4452;
12259: waveform_sig_loopback =3149;
12260: waveform_sig_loopback =4558;
12261: waveform_sig_loopback =4967;
12262: waveform_sig_loopback =3251;
12263: waveform_sig_loopback =3355;
12264: waveform_sig_loopback =5330;
12265: waveform_sig_loopback =4104;
12266: waveform_sig_loopback =2314;
12267: waveform_sig_loopback =4766;
12268: waveform_sig_loopback =4797;
12269: waveform_sig_loopback =2331;
12270: waveform_sig_loopback =6028;
12271: waveform_sig_loopback =1173;
12272: waveform_sig_loopback =2679;
12273: waveform_sig_loopback =6740;
12274: waveform_sig_loopback =2893;
12275: waveform_sig_loopback =2632;
12276: waveform_sig_loopback =2863;
12277: waveform_sig_loopback =4124;
12278: waveform_sig_loopback =4960;
12279: waveform_sig_loopback =2209;
12280: waveform_sig_loopback =2763;
12281: waveform_sig_loopback =4318;
12282: waveform_sig_loopback =2713;
12283: waveform_sig_loopback =3875;
12284: waveform_sig_loopback =2287;
12285: waveform_sig_loopback =3531;
12286: waveform_sig_loopback =3731;
12287: waveform_sig_loopback =2180;
12288: waveform_sig_loopback =3340;
12289: waveform_sig_loopback =3046;
12290: waveform_sig_loopback =2694;
12291: waveform_sig_loopback =2441;
12292: waveform_sig_loopback =4177;
12293: waveform_sig_loopback =1766;
12294: waveform_sig_loopback =2265;
12295: waveform_sig_loopback =3921;
12296: waveform_sig_loopback =2259;
12297: waveform_sig_loopback =2032;
12298: waveform_sig_loopback =3159;
12299: waveform_sig_loopback =2913;
12300: waveform_sig_loopback =1641;
12301: waveform_sig_loopback =2590;
12302: waveform_sig_loopback =3397;
12303: waveform_sig_loopback =1531;
12304: waveform_sig_loopback =1576;
12305: waveform_sig_loopback =3801;
12306: waveform_sig_loopback =2078;
12307: waveform_sig_loopback =697;
12308: waveform_sig_loopback =3328;
12309: waveform_sig_loopback =2633;
12310: waveform_sig_loopback =831;
12311: waveform_sig_loopback =4315;
12312: waveform_sig_loopback =-943;
12313: waveform_sig_loopback =1369;
12314: waveform_sig_loopback =4772;
12315: waveform_sig_loopback =1079;
12316: waveform_sig_loopback =1076;
12317: waveform_sig_loopback =788;
12318: waveform_sig_loopback =2540;
12319: waveform_sig_loopback =3276;
12320: waveform_sig_loopback =-6;
12321: waveform_sig_loopback =1275;
12322: waveform_sig_loopback =2369;
12323: waveform_sig_loopback =811;
12324: waveform_sig_loopback =2334;
12325: waveform_sig_loopback =42;
12326: waveform_sig_loopback =2051;
12327: waveform_sig_loopback =1912;
12328: waveform_sig_loopback =68;
12329: waveform_sig_loopback =1805;
12330: waveform_sig_loopback =1172;
12331: waveform_sig_loopback =910;
12332: waveform_sig_loopback =697;
12333: waveform_sig_loopback =2058;
12334: waveform_sig_loopback =68;
12335: waveform_sig_loopback =818;
12336: waveform_sig_loopback =1646;
12337: waveform_sig_loopback =455;
12338: waveform_sig_loopback =296;
12339: waveform_sig_loopback =1350;
12340: waveform_sig_loopback =1088;
12341: waveform_sig_loopback =-533;
12342: waveform_sig_loopback =977;
12343: waveform_sig_loopback =1655;
12344: waveform_sig_loopback =-641;
12345: waveform_sig_loopback =-217;
12346: waveform_sig_loopback =2133;
12347: waveform_sig_loopback =19;
12348: waveform_sig_loopback =-1128;
12349: waveform_sig_loopback =1513;
12350: waveform_sig_loopback =483;
12351: waveform_sig_loopback =-610;
12352: waveform_sig_loopback =2149;
12353: waveform_sig_loopback =-3007;
12354: waveform_sig_loopback =61;
12355: waveform_sig_loopback =2445;
12356: waveform_sig_loopback =-645;
12357: waveform_sig_loopback =-844;
12358: waveform_sig_loopback =-1274;
12359: waveform_sig_loopback =1121;
12360: waveform_sig_loopback =989;
12361: waveform_sig_loopback =-1924;
12362: waveform_sig_loopback =-219;
12363: waveform_sig_loopback =7;
12364: waveform_sig_loopback =-692;
12365: waveform_sig_loopback =285;
12366: waveform_sig_loopback =-1983;
12367: waveform_sig_loopback =593;
12368: waveform_sig_loopback =-464;
12369: waveform_sig_loopback =-1584;
12370: waveform_sig_loopback =-92;
12371: waveform_sig_loopback =-847;
12372: waveform_sig_loopback =-888;
12373: waveform_sig_loopback =-1255;
12374: waveform_sig_loopback =221;
12375: waveform_sig_loopback =-1952;
12376: waveform_sig_loopback =-929;
12377: waveform_sig_loopback =-450;
12378: waveform_sig_loopback =-1299;
12379: waveform_sig_loopback =-1668;
12380: waveform_sig_loopback =-730;
12381: waveform_sig_loopback =-547;
12382: waveform_sig_loopback =-2760;
12383: waveform_sig_loopback =-659;
12384: waveform_sig_loopback =-289;
12385: waveform_sig_loopback =-2893;
12386: waveform_sig_loopback =-1542;
12387: waveform_sig_loopback =-149;
12388: waveform_sig_loopback =-1962;
12389: waveform_sig_loopback =-2740;
12390: waveform_sig_loopback =-664;
12391: waveform_sig_loopback =-1137;
12392: waveform_sig_loopback =-2614;
12393: waveform_sig_loopback =94;
12394: waveform_sig_loopback =-4749;
12395: waveform_sig_loopback =-1884;
12396: waveform_sig_loopback =643;
12397: waveform_sig_loopback =-2621;
12398: waveform_sig_loopback =-2885;
12399: waveform_sig_loopback =-2885;
12400: waveform_sig_loopback =-845;
12401: waveform_sig_loopback =-957;
12402: waveform_sig_loopback =-3676;
12403: waveform_sig_loopback =-2090;
12404: waveform_sig_loopback =-1924;
12405: waveform_sig_loopback =-2390;
12406: waveform_sig_loopback =-1734;
12407: waveform_sig_loopback =-3796;
12408: waveform_sig_loopback =-1133;
12409: waveform_sig_loopback =-2537;
12410: waveform_sig_loopback =-3227;
12411: waveform_sig_loopback =-1946;
12412: waveform_sig_loopback =-2827;
12413: waveform_sig_loopback =-2556;
12414: waveform_sig_loopback =-3118;
12415: waveform_sig_loopback =-1697;
12416: waveform_sig_loopback =-3621;
12417: waveform_sig_loopback =-2951;
12418: waveform_sig_loopback =-2085;
12419: waveform_sig_loopback =-3139;
12420: waveform_sig_loopback =-3681;
12421: waveform_sig_loopback =-2049;
12422: waveform_sig_loopback =-2785;
12423: waveform_sig_loopback =-4498;
12424: waveform_sig_loopback =-2104;
12425: waveform_sig_loopback =-2520;
12426: waveform_sig_loopback =-4427;
12427: waveform_sig_loopback =-3272;
12428: waveform_sig_loopback =-2071;
12429: waveform_sig_loopback =-3522;
12430: waveform_sig_loopback =-4760;
12431: waveform_sig_loopback =-2213;
12432: waveform_sig_loopback =-2974;
12433: waveform_sig_loopback =-4484;
12434: waveform_sig_loopback =-1452;
12435: waveform_sig_loopback =-6789;
12436: waveform_sig_loopback =-3353;
12437: waveform_sig_loopback =-1129;
12438: waveform_sig_loopback =-4535;
12439: waveform_sig_loopback =-4605;
12440: waveform_sig_loopback =-4406;
12441: waveform_sig_loopback =-2597;
12442: waveform_sig_loopback =-2881;
12443: waveform_sig_loopback =-5290;
12444: waveform_sig_loopback =-3774;
12445: waveform_sig_loopback =-3596;
12446: waveform_sig_loopback =-4086;
12447: waveform_sig_loopback =-3661;
12448: waveform_sig_loopback =-5125;
12449: waveform_sig_loopback =-2899;
12450: waveform_sig_loopback =-4462;
12451: waveform_sig_loopback =-4582;
12452: waveform_sig_loopback =-3871;
12453: waveform_sig_loopback =-4297;
12454: waveform_sig_loopback =-4207;
12455: waveform_sig_loopback =-5039;
12456: waveform_sig_loopback =-2933;
12457: waveform_sig_loopback =-5566;
12458: waveform_sig_loopback =-4550;
12459: waveform_sig_loopback =-3449;
12460: waveform_sig_loopback =-5213;
12461: waveform_sig_loopback =-4925;
12462: waveform_sig_loopback =-3728;
12463: waveform_sig_loopback =-4615;
12464: waveform_sig_loopback =-5695;
12465: waveform_sig_loopback =-3957;
12466: waveform_sig_loopback =-4008;
12467: waveform_sig_loopback =-6029;
12468: waveform_sig_loopback =-4879;
12469: waveform_sig_loopback =-3491;
12470: waveform_sig_loopback =-5271;
12471: waveform_sig_loopback =-6232;
12472: waveform_sig_loopback =-3568;
12473: waveform_sig_loopback =-4659;
12474: waveform_sig_loopback =-5915;
12475: waveform_sig_loopback =-2996;
12476: waveform_sig_loopback =-8360;
12477: waveform_sig_loopback =-4682;
12478: waveform_sig_loopback =-2590;
12479: waveform_sig_loopback =-6148;
12480: waveform_sig_loopback =-6112;
12481: waveform_sig_loopback =-5679;
12482: waveform_sig_loopback =-4222;
12483: waveform_sig_loopback =-4192;
12484: waveform_sig_loopback =-6826;
12485: waveform_sig_loopback =-5365;
12486: waveform_sig_loopback =-4738;
12487: waveform_sig_loopback =-5763;
12488: waveform_sig_loopback =-5008;
12489: waveform_sig_loopback =-6411;
12490: waveform_sig_loopback =-4644;
12491: waveform_sig_loopback =-5450;
12492: waveform_sig_loopback =-6103;
12493: waveform_sig_loopback =-5400;
12494: waveform_sig_loopback =-5279;
12495: waveform_sig_loopback =-6107;
12496: waveform_sig_loopback =-5921;
12497: waveform_sig_loopback =-4429;
12498: waveform_sig_loopback =-7156;
12499: waveform_sig_loopback =-5409;
12500: waveform_sig_loopback =-5183;
12501: waveform_sig_loopback =-6367;
12502: waveform_sig_loopback =-6237;
12503: waveform_sig_loopback =-5083;
12504: waveform_sig_loopback =-5889;
12505: waveform_sig_loopback =-7072;
12506: waveform_sig_loopback =-5084;
12507: waveform_sig_loopback =-5437;
12508: waveform_sig_loopback =-7187;
12509: waveform_sig_loopback =-6171;
12510: waveform_sig_loopback =-4639;
12511: waveform_sig_loopback =-6527;
12512: waveform_sig_loopback =-7637;
12513: waveform_sig_loopback =-4385;
12514: waveform_sig_loopback =-6247;
12515: waveform_sig_loopback =-6921;
12516: waveform_sig_loopback =-4032;
12517: waveform_sig_loopback =-10074;
12518: waveform_sig_loopback =-5182;
12519: waveform_sig_loopback =-3976;
12520: waveform_sig_loopback =-7583;
12521: waveform_sig_loopback =-6812;
12522: waveform_sig_loopback =-7145;
12523: waveform_sig_loopback =-5075;
12524: waveform_sig_loopback =-5255;
12525: waveform_sig_loopback =-8356;
12526: waveform_sig_loopback =-5855;
12527: waveform_sig_loopback =-6110;
12528: waveform_sig_loopback =-6853;
12529: waveform_sig_loopback =-5799;
12530: waveform_sig_loopback =-7751;
12531: waveform_sig_loopback =-5409;
12532: waveform_sig_loopback =-6603;
12533: waveform_sig_loopback =-7289;
12534: waveform_sig_loopback =-6094;
12535: waveform_sig_loopback =-6508;
12536: waveform_sig_loopback =-7050;
12537: waveform_sig_loopback =-6728;
12538: waveform_sig_loopback =-5562;
12539: waveform_sig_loopback =-8042;
12540: waveform_sig_loopback =-6226;
12541: waveform_sig_loopback =-6175;
12542: waveform_sig_loopback =-7287;
12543: waveform_sig_loopback =-6958;
12544: waveform_sig_loopback =-6140;
12545: waveform_sig_loopback =-6703;
12546: waveform_sig_loopback =-7853;
12547: waveform_sig_loopback =-6056;
12548: waveform_sig_loopback =-6097;
12549: waveform_sig_loopback =-8216;
12550: waveform_sig_loopback =-6845;
12551: waveform_sig_loopback =-5357;
12552: waveform_sig_loopback =-7673;
12553: waveform_sig_loopback =-8116;
12554: waveform_sig_loopback =-5100;
12555: waveform_sig_loopback =-7421;
12556: waveform_sig_loopback =-7203;
12557: waveform_sig_loopback =-5153;
12558: waveform_sig_loopback =-10864;
12559: waveform_sig_loopback =-5421;
12560: waveform_sig_loopback =-5263;
12561: waveform_sig_loopback =-7911;
12562: waveform_sig_loopback =-7595;
12563: waveform_sig_loopback =-8027;
12564: waveform_sig_loopback =-5268;
12565: waveform_sig_loopback =-6375;
12566: waveform_sig_loopback =-8863;
12567: waveform_sig_loopback =-6303;
12568: waveform_sig_loopback =-7122;
12569: waveform_sig_loopback =-7075;
12570: waveform_sig_loopback =-6668;
12571: waveform_sig_loopback =-8411;
12572: waveform_sig_loopback =-5684;
12573: waveform_sig_loopback =-7511;
12574: waveform_sig_loopback =-7640;
12575: waveform_sig_loopback =-6683;
12576: waveform_sig_loopback =-7076;
12577: waveform_sig_loopback =-7558;
12578: waveform_sig_loopback =-7110;
12579: waveform_sig_loopback =-6205;
12580: waveform_sig_loopback =-8564;
12581: waveform_sig_loopback =-6419;
12582: waveform_sig_loopback =-6913;
12583: waveform_sig_loopback =-7560;
12584: waveform_sig_loopback =-7476;
12585: waveform_sig_loopback =-6615;
12586: waveform_sig_loopback =-6787;
12587: waveform_sig_loopback =-8682;
12588: waveform_sig_loopback =-6122;
12589: waveform_sig_loopback =-6549;
12590: waveform_sig_loopback =-8860;
12591: waveform_sig_loopback =-6726;
12592: waveform_sig_loopback =-6026;
12593: waveform_sig_loopback =-8043;
12594: waveform_sig_loopback =-8139;
12595: waveform_sig_loopback =-5695;
12596: waveform_sig_loopback =-7602;
12597: waveform_sig_loopback =-7303;
12598: waveform_sig_loopback =-5822;
12599: waveform_sig_loopback =-10802;
12600: waveform_sig_loopback =-5643;
12601: waveform_sig_loopback =-5622;
12602: waveform_sig_loopback =-7929;
12603: waveform_sig_loopback =-8152;
12604: waveform_sig_loopback =-7932;
12605: waveform_sig_loopback =-5408;
12606: waveform_sig_loopback =-6802;
12607: waveform_sig_loopback =-8837;
12608: waveform_sig_loopback =-6502;
12609: waveform_sig_loopback =-7384;
12610: waveform_sig_loopback =-6916;
12611: waveform_sig_loopback =-7029;
12612: waveform_sig_loopback =-8437;
12613: waveform_sig_loopback =-5616;
12614: waveform_sig_loopback =-7857;
12615: waveform_sig_loopback =-7503;
12616: waveform_sig_loopback =-6724;
12617: waveform_sig_loopback =-7320;
12618: waveform_sig_loopback =-7386;
12619: waveform_sig_loopback =-7186;
12620: waveform_sig_loopback =-6392;
12621: waveform_sig_loopback =-8247;
12622: waveform_sig_loopback =-6751;
12623: waveform_sig_loopback =-6758;
12624: waveform_sig_loopback =-7416;
12625: waveform_sig_loopback =-7685;
12626: waveform_sig_loopback =-6121;
12627: waveform_sig_loopback =-7167;
12628: waveform_sig_loopback =-8452;
12629: waveform_sig_loopback =-5760;
12630: waveform_sig_loopback =-6818;
12631: waveform_sig_loopback =-8612;
12632: waveform_sig_loopback =-6514;
12633: waveform_sig_loopback =-6097;
12634: waveform_sig_loopback =-7825;
12635: waveform_sig_loopback =-7952;
12636: waveform_sig_loopback =-5679;
12637: waveform_sig_loopback =-7268;
12638: waveform_sig_loopback =-7260;
12639: waveform_sig_loopback =-5903;
12640: waveform_sig_loopback =-10278;
12641: waveform_sig_loopback =-5547;
12642: waveform_sig_loopback =-5354;
12643: waveform_sig_loopback =-7987;
12644: waveform_sig_loopback =-7960;
12645: waveform_sig_loopback =-7125;
12646: waveform_sig_loopback =-5541;
12647: waveform_sig_loopback =-6674;
12648: waveform_sig_loopback =-8238;
12649: waveform_sig_loopback =-6284;
12650: waveform_sig_loopback =-6987;
12651: waveform_sig_loopback =-6679;
12652: waveform_sig_loopback =-6796;
12653: waveform_sig_loopback =-7710;
12654: waveform_sig_loopback =-5484;
12655: waveform_sig_loopback =-7558;
12656: waveform_sig_loopback =-6830;
12657: waveform_sig_loopback =-6480;
12658: waveform_sig_loopback =-6888;
12659: waveform_sig_loopback =-6959;
12660: waveform_sig_loopback =-6727;
12661: waveform_sig_loopback =-5865;
12662: waveform_sig_loopback =-7798;
12663: waveform_sig_loopback =-6436;
12664: waveform_sig_loopback =-5954;
12665: waveform_sig_loopback =-7133;
12666: waveform_sig_loopback =-7223;
12667: waveform_sig_loopback =-5297;
12668: waveform_sig_loopback =-7144;
12669: waveform_sig_loopback =-7472;
12670: waveform_sig_loopback =-5264;
12671: waveform_sig_loopback =-6545;
12672: waveform_sig_loopback =-7582;
12673: waveform_sig_loopback =-6186;
12674: waveform_sig_loopback =-5361;
12675: waveform_sig_loopback =-7148;
12676: waveform_sig_loopback =-7498;
12677: waveform_sig_loopback =-4632;
12678: waveform_sig_loopback =-6910;
12679: waveform_sig_loopback =-6384;
12680: waveform_sig_loopback =-4997;
12681: waveform_sig_loopback =-9913;
12682: waveform_sig_loopback =-4563;
12683: waveform_sig_loopback =-4539;
12684: waveform_sig_loopback =-7320;
12685: waveform_sig_loopback =-7187;
12686: waveform_sig_loopback =-6386;
12687: waveform_sig_loopback =-4798;
12688: waveform_sig_loopback =-5642;
12689: waveform_sig_loopback =-7695;
12690: waveform_sig_loopback =-5543;
12691: waveform_sig_loopback =-5938;
12692: waveform_sig_loopback =-5986;
12693: waveform_sig_loopback =-6001;
12694: waveform_sig_loopback =-6767;
12695: waveform_sig_loopback =-4753;
12696: waveform_sig_loopback =-6543;
12697: waveform_sig_loopback =-6010;
12698: waveform_sig_loopback =-5776;
12699: waveform_sig_loopback =-5681;
12700: waveform_sig_loopback =-6211;
12701: waveform_sig_loopback =-5875;
12702: waveform_sig_loopback =-4762;
12703: waveform_sig_loopback =-7130;
12704: waveform_sig_loopback =-5246;
12705: waveform_sig_loopback =-5025;
12706: waveform_sig_loopback =-6530;
12707: waveform_sig_loopback =-5698;
12708: waveform_sig_loopback =-4610;
12709: waveform_sig_loopback =-6252;
12710: waveform_sig_loopback =-6055;
12711: waveform_sig_loopback =-4626;
12712: waveform_sig_loopback =-5314;
12713: waveform_sig_loopback =-6609;
12714: waveform_sig_loopback =-5203;
12715: waveform_sig_loopback =-4002;
12716: waveform_sig_loopback =-6482;
12717: waveform_sig_loopback =-6238;
12718: waveform_sig_loopback =-3355;
12719: waveform_sig_loopback =-6207;
12720: waveform_sig_loopback =-4868;
12721: waveform_sig_loopback =-4131;
12722: waveform_sig_loopback =-8818;
12723: waveform_sig_loopback =-3036;
12724: waveform_sig_loopback =-3713;
12725: waveform_sig_loopback =-6167;
12726: waveform_sig_loopback =-5882;
12727: waveform_sig_loopback =-5317;
12728: waveform_sig_loopback =-3502;
12729: waveform_sig_loopback =-4399;
12730: waveform_sig_loopback =-6652;
12731: waveform_sig_loopback =-4147;
12732: waveform_sig_loopback =-4765;
12733: waveform_sig_loopback =-4804;
12734: waveform_sig_loopback =-4673;
12735: waveform_sig_loopback =-5587;
12736: waveform_sig_loopback =-3472;
12737: waveform_sig_loopback =-5166;
12738: waveform_sig_loopback =-4867;
12739: waveform_sig_loopback =-4454;
12740: waveform_sig_loopback =-4176;
12741: waveform_sig_loopback =-5285;
12742: waveform_sig_loopback =-4098;
12743: waveform_sig_loopback =-3650;
12744: waveform_sig_loopback =-5988;
12745: waveform_sig_loopback =-3301;
12746: waveform_sig_loopback =-4245;
12747: waveform_sig_loopback =-4863;
12748: waveform_sig_loopback =-4254;
12749: waveform_sig_loopback =-3529;
12750: waveform_sig_loopback =-4401;
12751: waveform_sig_loopback =-5091;
12752: waveform_sig_loopback =-2982;
12753: waveform_sig_loopback =-3790;
12754: waveform_sig_loopback =-5530;
12755: waveform_sig_loopback =-3381;
12756: waveform_sig_loopback =-2762;
12757: waveform_sig_loopback =-5100;
12758: waveform_sig_loopback =-4598;
12759: waveform_sig_loopback =-2013;
12760: waveform_sig_loopback =-4783;
12761: waveform_sig_loopback =-3229;
12762: waveform_sig_loopback =-2933;
12763: waveform_sig_loopback =-7363;
12764: waveform_sig_loopback =-1199;
12765: waveform_sig_loopback =-2508;
12766: waveform_sig_loopback =-4664;
12767: waveform_sig_loopback =-4161;
12768: waveform_sig_loopback =-4012;
12769: waveform_sig_loopback =-1645;
12770: waveform_sig_loopback =-3100;
12771: waveform_sig_loopback =-5309;
12772: waveform_sig_loopback =-2082;
12773: waveform_sig_loopback =-3696;
12774: waveform_sig_loopback =-2921;
12775: waveform_sig_loopback =-3046;
12776: waveform_sig_loopback =-4326;
12777: waveform_sig_loopback =-1418;
12778: waveform_sig_loopback =-3915;
12779: waveform_sig_loopback =-3234;
12780: waveform_sig_loopback =-2517;
12781: waveform_sig_loopback =-3040;
12782: waveform_sig_loopback =-3319;
12783: waveform_sig_loopback =-2382;
12784: waveform_sig_loopback =-2414;
12785: waveform_sig_loopback =-3911;
12786: waveform_sig_loopback =-1960;
12787: waveform_sig_loopback =-2472;
12788: waveform_sig_loopback =-3074;
12789: waveform_sig_loopback =-2905;
12790: waveform_sig_loopback =-1632;
12791: waveform_sig_loopback =-2882;
12792: waveform_sig_loopback =-3351;
12793: waveform_sig_loopback =-1168;
12794: waveform_sig_loopback =-2306;
12795: waveform_sig_loopback =-3831;
12796: waveform_sig_loopback =-1454;
12797: waveform_sig_loopback =-1185;
12798: waveform_sig_loopback =-3519;
12799: waveform_sig_loopback =-2613;
12800: waveform_sig_loopback =-456;
12801: waveform_sig_loopback =-3101;
12802: waveform_sig_loopback =-1097;
12803: waveform_sig_loopback =-1750;
12804: waveform_sig_loopback =-5227;
12805: waveform_sig_loopback =595;
12806: waveform_sig_loopback =-1043;
12807: waveform_sig_loopback =-2536;
12808: waveform_sig_loopback =-2925;
12809: waveform_sig_loopback =-1973;
12810: waveform_sig_loopback =296;
12811: waveform_sig_loopback =-1862;
12812: waveform_sig_loopback =-3013;
12813: waveform_sig_loopback =-532;
12814: waveform_sig_loopback =-2013;
12815: waveform_sig_loopback =-708;
12816: waveform_sig_loopback =-1853;
12817: waveform_sig_loopback =-2121;
12818: waveform_sig_loopback =425;
12819: waveform_sig_loopback =-2542;
12820: waveform_sig_loopback =-922;
12821: waveform_sig_loopback =-1049;
12822: waveform_sig_loopback =-1130;
12823: waveform_sig_loopback =-1442;
12824: waveform_sig_loopback =-806;
12825: waveform_sig_loopback =-385;
12826: waveform_sig_loopback =-2095;
12827: waveform_sig_loopback =-173;
12828: waveform_sig_loopback =-553;
12829: waveform_sig_loopback =-1360;
12830: waveform_sig_loopback =-950;
12831: waveform_sig_loopback =355;
12832: waveform_sig_loopback =-1278;
12833: waveform_sig_loopback =-1528;
12834: waveform_sig_loopback =861;
12835: waveform_sig_loopback =-649;
12836: waveform_sig_loopback =-1977;
12837: waveform_sig_loopback =572;
12838: waveform_sig_loopback =407;
12839: waveform_sig_loopback =-1492;
12840: waveform_sig_loopback =-669;
12841: waveform_sig_loopback =1190;
12842: waveform_sig_loopback =-984;
12843: waveform_sig_loopback =561;
12844: waveform_sig_loopback =36;
12845: waveform_sig_loopback =-3054;
12846: waveform_sig_loopback =2200;
12847: waveform_sig_loopback =1086;
12848: waveform_sig_loopback =-826;
12849: waveform_sig_loopback =-1116;
12850: waveform_sig_loopback =388;
12851: waveform_sig_loopback =1739;
12852: waveform_sig_loopback =200;
12853: waveform_sig_loopback =-1017;
12854: waveform_sig_loopback =1049;
12855: waveform_sig_loopback =209;
12856: waveform_sig_loopback =956;
12857: waveform_sig_loopback =6;
12858: waveform_sig_loopback =79;
12859: waveform_sig_loopback =1939;
12860: waveform_sig_loopback =-385;
12861: waveform_sig_loopback =917;
12862: waveform_sig_loopback =775;
12863: waveform_sig_loopback =879;
12864: waveform_sig_loopback =368;
12865: waveform_sig_loopback =1236;
12866: waveform_sig_loopback =1356;
12867: waveform_sig_loopback =-149;
12868: waveform_sig_loopback =1620;
12869: waveform_sig_loopback =1447;
12870: waveform_sig_loopback =392;
12871: waveform_sig_loopback =890;
12872: waveform_sig_loopback =2476;
12873: waveform_sig_loopback =216;
12874: waveform_sig_loopback =735;
12875: waveform_sig_loopback =2708;
12876: waveform_sig_loopback =881;
12877: waveform_sig_loopback =418;
12878: waveform_sig_loopback =2123;
12879: waveform_sig_loopback =2364;
12880: waveform_sig_loopback =507;
12881: waveform_sig_loopback =939;
12882: waveform_sig_loopback =3463;
12883: waveform_sig_loopback =531;
12884: waveform_sig_loopback =2553;
12885: waveform_sig_loopback =2004;
12886: waveform_sig_loopback =-1478;
12887: waveform_sig_loopback =4483;
12888: waveform_sig_loopback =2763;
12889: waveform_sig_loopback =782;
12890: waveform_sig_loopback =1110;
12891: waveform_sig_loopback =2106;
12892: waveform_sig_loopback =3599;
12893: waveform_sig_loopback =2050;
12894: waveform_sig_loopback =781;
12895: waveform_sig_loopback =3030;
12896: waveform_sig_loopback =2024;
12897: waveform_sig_loopback =2690;
12898: waveform_sig_loopback =1899;
12899: waveform_sig_loopback =2049;
12900: waveform_sig_loopback =3556;
12901: waveform_sig_loopback =1577;
12902: waveform_sig_loopback =2745;
12903: waveform_sig_loopback =2510;
12904: waveform_sig_loopback =2962;
12905: waveform_sig_loopback =1923;
12906: waveform_sig_loopback =3176;
12907: waveform_sig_loopback =3291;
12908: waveform_sig_loopback =1406;
12909: waveform_sig_loopback =3778;
12910: waveform_sig_loopback =3061;
12911: waveform_sig_loopback =2081;
12912: waveform_sig_loopback =3163;
12913: waveform_sig_loopback =3856;
12914: waveform_sig_loopback =2187;
12915: waveform_sig_loopback =2701;
12916: waveform_sig_loopback =4282;
12917: waveform_sig_loopback =2886;
12918: waveform_sig_loopback =2076;
12919: waveform_sig_loopback =4001;
12920: waveform_sig_loopback =4231;
12921: waveform_sig_loopback =2016;
12922: waveform_sig_loopback =2882;
12923: waveform_sig_loopback =5363;
12924: waveform_sig_loopback =1964;
12925: waveform_sig_loopback =4637;
12926: waveform_sig_loopback =3439;
12927: waveform_sig_loopback =286;
12928: waveform_sig_loopback =6645;
12929: waveform_sig_loopback =4056;
12930: waveform_sig_loopback =2602;
12931: waveform_sig_loopback =3019;
12932: waveform_sig_loopback =3716;
12933: waveform_sig_loopback =5442;
12934: waveform_sig_loopback =3575;
12935: waveform_sig_loopback =2465;
12936: waveform_sig_loopback =4981;
12937: waveform_sig_loopback =3605;
12938: waveform_sig_loopback =4370;
12939: waveform_sig_loopback =3688;
12940: waveform_sig_loopback =3760;
12941: waveform_sig_loopback =5148;
12942: waveform_sig_loopback =3430;
12943: waveform_sig_loopback =4208;
12944: waveform_sig_loopback =4360;
12945: waveform_sig_loopback =4620;
12946: waveform_sig_loopback =3292;
12947: waveform_sig_loopback =5356;
12948: waveform_sig_loopback =4471;
12949: waveform_sig_loopback =3130;
12950: waveform_sig_loopback =5669;
12951: waveform_sig_loopback =4308;
12952: waveform_sig_loopback =4057;
12953: waveform_sig_loopback =4601;
12954: waveform_sig_loopback =5424;
12955: waveform_sig_loopback =3962;
12956: waveform_sig_loopback =4095;
12957: waveform_sig_loopback =6018;
12958: waveform_sig_loopback =4344;
12959: waveform_sig_loopback =3593;
12960: waveform_sig_loopback =5776;
12961: waveform_sig_loopback =5657;
12962: waveform_sig_loopback =3516;
12963: waveform_sig_loopback =4658;
12964: waveform_sig_loopback =6874;
12965: waveform_sig_loopback =3318;
12966: waveform_sig_loopback =6563;
12967: waveform_sig_loopback =4586;
12968: waveform_sig_loopback =1918;
12969: waveform_sig_loopback =8436;
12970: waveform_sig_loopback =5164;
12971: waveform_sig_loopback =4281;
12972: waveform_sig_loopback =4462;
12973: waveform_sig_loopback =5041;
12974: waveform_sig_loopback =7269;
12975: waveform_sig_loopback =4697;
12976: waveform_sig_loopback =4003;
12977: waveform_sig_loopback =6579;
12978: waveform_sig_loopback =4697;
12979: waveform_sig_loopback =6097;
12980: waveform_sig_loopback =4949;
12981: waveform_sig_loopback =5010;
12982: waveform_sig_loopback =6874;
12983: waveform_sig_loopback =4455;
12984: waveform_sig_loopback =5673;
12985: waveform_sig_loopback =5881;
12986: waveform_sig_loopback =5627;
12987: waveform_sig_loopback =4994;
12988: waveform_sig_loopback =6473;
12989: waveform_sig_loopback =5556;
12990: waveform_sig_loopback =4924;
12991: waveform_sig_loopback =6762;
12992: waveform_sig_loopback =5520;
12993: waveform_sig_loopback =5189;
12994: waveform_sig_loopback =6082;
12995: waveform_sig_loopback =6756;
12996: waveform_sig_loopback =5027;
12997: waveform_sig_loopback =5289;
12998: waveform_sig_loopback =7430;
12999: waveform_sig_loopback =5663;
13000: waveform_sig_loopback =4534;
13001: waveform_sig_loopback =7226;
13002: waveform_sig_loopback =6755;
13003: waveform_sig_loopback =4640;
13004: waveform_sig_loopback =6155;
13005: waveform_sig_loopback =7566;
13006: waveform_sig_loopback =4798;
13007: waveform_sig_loopback =7918;
13008: waveform_sig_loopback =5132;
13009: waveform_sig_loopback =3690;
13010: waveform_sig_loopback =9369;
13011: waveform_sig_loopback =6201;
13012: waveform_sig_loopback =5648;
13013: waveform_sig_loopback =5119;
13014: waveform_sig_loopback =6675;
13015: waveform_sig_loopback =8315;
13016: waveform_sig_loopback =5428;
13017: waveform_sig_loopback =5498;
13018: waveform_sig_loopback =7373;
13019: waveform_sig_loopback =5862;
13020: waveform_sig_loopback =7267;
13021: waveform_sig_loopback =5578;
13022: waveform_sig_loopback =6452;
13023: waveform_sig_loopback =7801;
13024: waveform_sig_loopback =5302;
13025: waveform_sig_loopback =6928;
13026: waveform_sig_loopback =6669;
13027: waveform_sig_loopback =6592;
13028: waveform_sig_loopback =6002;
13029: waveform_sig_loopback =7494;
13030: waveform_sig_loopback =6488;
13031: waveform_sig_loopback =5890;
13032: waveform_sig_loopback =7484;
13033: waveform_sig_loopback =6633;
13034: waveform_sig_loopback =6257;
13035: waveform_sig_loopback =6587;
13036: waveform_sig_loopback =7876;
13037: waveform_sig_loopback =5709;
13038: waveform_sig_loopback =6375;
13039: waveform_sig_loopback =8369;
13040: waveform_sig_loopback =5991;
13041: waveform_sig_loopback =5839;
13042: waveform_sig_loopback =8065;
13043: waveform_sig_loopback =7254;
13044: waveform_sig_loopback =5594;
13045: waveform_sig_loopback =6997;
13046: waveform_sig_loopback =8313;
13047: waveform_sig_loopback =5608;
13048: waveform_sig_loopback =8533;
13049: waveform_sig_loopback =5818;
13050: waveform_sig_loopback =4688;
13051: waveform_sig_loopback =9821;
13052: waveform_sig_loopback =7168;
13053: waveform_sig_loopback =6214;
13054: waveform_sig_loopback =5752;
13055: waveform_sig_loopback =7609;
13056: waveform_sig_loopback =8631;
13057: waveform_sig_loopback =6235;
13058: waveform_sig_loopback =6252;
13059: waveform_sig_loopback =7759;
13060: waveform_sig_loopback =6690;
13061: waveform_sig_loopback =7868;
13062: waveform_sig_loopback =6096;
13063: waveform_sig_loopback =7260;
13064: waveform_sig_loopback =8063;
13065: waveform_sig_loopback =6033;
13066: waveform_sig_loopback =7622;
13067: waveform_sig_loopback =6981;
13068: waveform_sig_loopback =7285;
13069: waveform_sig_loopback =6557;
13070: waveform_sig_loopback =7988;
13071: waveform_sig_loopback =6982;
13072: waveform_sig_loopback =6397;
13073: waveform_sig_loopback =7956;
13074: waveform_sig_loopback =7324;
13075: waveform_sig_loopback =6447;
13076: waveform_sig_loopback =7263;
13077: waveform_sig_loopback =8371;
13078: waveform_sig_loopback =5838;
13079: waveform_sig_loopback =7111;
13080: waveform_sig_loopback =8557;
13081: waveform_sig_loopback =6258;
13082: waveform_sig_loopback =6561;
13083: waveform_sig_loopback =8106;
13084: waveform_sig_loopback =7708;
13085: waveform_sig_loopback =5978;
13086: waveform_sig_loopback =7157;
13087: waveform_sig_loopback =8873;
13088: waveform_sig_loopback =5677;
13089: waveform_sig_loopback =8986;
13090: waveform_sig_loopback =5984;
13091: waveform_sig_loopback =4937;
13092: waveform_sig_loopback =10291;
13093: waveform_sig_loopback =7230;
13094: waveform_sig_loopback =6215;
13095: waveform_sig_loopback =6237;
13096: waveform_sig_loopback =7858;
13097: waveform_sig_loopback =8594;
13098: waveform_sig_loopback =6546;
13099: waveform_sig_loopback =6303;
13100: waveform_sig_loopback =8007;
13101: waveform_sig_loopback =6933;
13102: waveform_sig_loopback =7652;
13103: waveform_sig_loopback =6473;
13104: waveform_sig_loopback =7390;
13105: waveform_sig_loopback =7906;
13106: waveform_sig_loopback =6253;
13107: waveform_sig_loopback =7641;
13108: waveform_sig_loopback =7069;
13109: waveform_sig_loopback =7296;
13110: waveform_sig_loopback =6496;
13111: waveform_sig_loopback =8092;
13112: waveform_sig_loopback =7072;
13113: waveform_sig_loopback =6118;
13114: waveform_sig_loopback =8152;
13115: waveform_sig_loopback =7147;
13116: waveform_sig_loopback =6313;
13117: waveform_sig_loopback =7584;
13118: waveform_sig_loopback =7928;
13119: waveform_sig_loopback =5820;
13120: waveform_sig_loopback =7286;
13121: waveform_sig_loopback =8292;
13122: waveform_sig_loopback =6184;
13123: waveform_sig_loopback =6409;
13124: waveform_sig_loopback =8103;
13125: waveform_sig_loopback =7585;
13126: waveform_sig_loopback =5651;
13127: waveform_sig_loopback =7137;
13128: waveform_sig_loopback =8814;
13129: waveform_sig_loopback =5228;
13130: waveform_sig_loopback =8941;
13131: waveform_sig_loopback =5725;
13132: waveform_sig_loopback =4732;
13133: waveform_sig_loopback =10134;
13134: waveform_sig_loopback =6812;
13135: waveform_sig_loopback =5928;
13136: waveform_sig_loopback =6171;
13137: waveform_sig_loopback =7226;
13138: waveform_sig_loopback =8515;
13139: waveform_sig_loopback =6167;
13140: waveform_sig_loopback =5821;
13141: waveform_sig_loopback =7917;
13142: waveform_sig_loopback =6420;
13143: waveform_sig_loopback =7380;
13144: waveform_sig_loopback =6011;
13145: waveform_sig_loopback =7054;
13146: waveform_sig_loopback =7498;
13147: waveform_sig_loopback =5879;
13148: waveform_sig_loopback =7147;
13149: waveform_sig_loopback =6629;
13150: waveform_sig_loopback =7036;
13151: waveform_sig_loopback =5856;
13152: waveform_sig_loopback =7800;
13153: waveform_sig_loopback =6409;
13154: waveform_sig_loopback =5710;
13155: waveform_sig_loopback =7993;
13156: waveform_sig_loopback =6251;
13157: waveform_sig_loopback =5853;
13158: waveform_sig_loopback =7397;
13159: waveform_sig_loopback =6972;
13160: waveform_sig_loopback =5519;
13161: waveform_sig_loopback =6719;
13162: waveform_sig_loopback =7598;
13163: waveform_sig_loopback =5906;
13164: waveform_sig_loopback =5398;
13165: waveform_sig_loopback =7822;
13166: waveform_sig_loopback =6945;
13167: waveform_sig_loopback =4642;
13168: waveform_sig_loopback =6992;
13169: waveform_sig_loopback =7725;
13170: waveform_sig_loopback =4696;
13171: waveform_sig_loopback =8443;
13172: waveform_sig_loopback =4412;
13173: waveform_sig_loopback =4532;
13174: waveform_sig_loopback =9469;
13175: waveform_sig_loopback =5789;
13176: waveform_sig_loopback =5372;
13177: waveform_sig_loopback =5373;
13178: waveform_sig_loopback =6600;
13179: waveform_sig_loopback =7878;
13180: waveform_sig_loopback =5105;
13181: waveform_sig_loopback =5173;
13182: waveform_sig_loopback =7205;
13183: waveform_sig_loopback =5455;
13184: waveform_sig_loopback =6668;
13185: waveform_sig_loopback =5178;
13186: waveform_sig_loopback =6149;
13187: waveform_sig_loopback =6777;
13188: waveform_sig_loopback =5009;
13189: waveform_sig_loopback =6158;
13190: waveform_sig_loopback =6032;
13191: waveform_sig_loopback =5867;
13192: waveform_sig_loopback =4999;
13193: waveform_sig_loopback =7210;
13194: waveform_sig_loopback =4913;
13195: waveform_sig_loopback =5203;
13196: waveform_sig_loopback =6912;
13197: waveform_sig_loopback =5080;
13198: waveform_sig_loopback =5284;
13199: waveform_sig_loopback =5955;
13200: waveform_sig_loopback =6179;
13201: waveform_sig_loopback =4607;
13202: waveform_sig_loopback =5399;
13203: waveform_sig_loopback =6864;
13204: waveform_sig_loopback =4611;
13205: waveform_sig_loopback =4391;
13206: waveform_sig_loopback =7022;
13207: waveform_sig_loopback =5492;
13208: waveform_sig_loopback =3748;
13209: waveform_sig_loopback =6101;
13210: waveform_sig_loopback =6312;
13211: waveform_sig_loopback =3849;
13212: waveform_sig_loopback =7313;
13213: waveform_sig_loopback =3063;
13214: waveform_sig_loopback =3751;
13215: waveform_sig_loopback =8184;
13216: waveform_sig_loopback =4621;
13217: waveform_sig_loopback =4285;
13218: waveform_sig_loopback =4116;
13219: waveform_sig_loopback =5462;
13220: waveform_sig_loopback =6827;
13221: waveform_sig_loopback =3620;
13222: waveform_sig_loopback =4186;
13223: waveform_sig_loopback =6016;
13224: waveform_sig_loopback =3937;
13225: waveform_sig_loopback =5846;
13226: waveform_sig_loopback =3577;
13227: waveform_sig_loopback =5000;
13228: waveform_sig_loopback =5744;
13229: waveform_sig_loopback =3293;
13230: waveform_sig_loopback =5258;
13231: waveform_sig_loopback =4615;
13232: waveform_sig_loopback =4292;
13233: waveform_sig_loopback =4212;
13234: waveform_sig_loopback =5449;
13235: waveform_sig_loopback =3698;
13236: waveform_sig_loopback =4137;
13237: waveform_sig_loopback =5095;
13238: waveform_sig_loopback =4149;
13239: waveform_sig_loopback =3679;
13240: waveform_sig_loopback =4625;
13241: waveform_sig_loopback =5014;
13242: waveform_sig_loopback =2839;
13243: waveform_sig_loopback =4367;
13244: waveform_sig_loopback =5385;
13245: waveform_sig_loopback =3010;
13246: waveform_sig_loopback =3207;
13247: waveform_sig_loopback =5512;
13248: waveform_sig_loopback =3984;
13249: waveform_sig_loopback =2304;
13250: waveform_sig_loopback =4762;
13251: waveform_sig_loopback =4640;
13252: waveform_sig_loopback =2541;
13253: waveform_sig_loopback =5853;
13254: waveform_sig_loopback =1172;
13255: waveform_sig_loopback =2848;
13256: waveform_sig_loopback =6387;
13257: waveform_sig_loopback =3053;
13258: waveform_sig_loopback =2985;
13259: waveform_sig_loopback =2242;
13260: waveform_sig_loopback =4456;
13261: waveform_sig_loopback =4957;
13262: waveform_sig_loopback =1850;
13263: waveform_sig_loopback =3197;
13264: waveform_sig_loopback =3875;
13265: waveform_sig_loopback =2768;
13266: waveform_sig_loopback =4170;
13267: waveform_sig_loopback =1685;
13268: waveform_sig_loopback =4085;
13269: waveform_sig_loopback =3563;
13270: waveform_sig_loopback =1876;
13271: waveform_sig_loopback =3875;
13272: waveform_sig_loopback =2641;
13273: waveform_sig_loopback =3050;
13274: waveform_sig_loopback =2345;
13275: waveform_sig_loopback =3810;
13276: waveform_sig_loopback =2217;
13277: waveform_sig_loopback =2254;
13278: waveform_sig_loopback =3631;
13279: waveform_sig_loopback =2351;
13280: waveform_sig_loopback =2042;
13281: waveform_sig_loopback =3080;
13282: waveform_sig_loopback =3220;
13283: waveform_sig_loopback =1175;
13284: waveform_sig_loopback =2674;
13285: waveform_sig_loopback =3759;
13286: waveform_sig_loopback =1088;
13287: waveform_sig_loopback =1793;
13288: waveform_sig_loopback =3846;
13289: waveform_sig_loopback =1918;
13290: waveform_sig_loopback =1011;
13291: waveform_sig_loopback =2910;
13292: waveform_sig_loopback =2888;
13293: waveform_sig_loopback =1065;
13294: waveform_sig_loopback =3748;
13295: waveform_sig_loopback =-292;
13296: waveform_sig_loopback =1120;
13297: waveform_sig_loopback =4478;
13298: waveform_sig_loopback =1643;
13299: waveform_sig_loopback =745;
13300: waveform_sig_loopback =844;
13301: waveform_sig_loopback =2802;
13302: waveform_sig_loopback =2837;
13303: waveform_sig_loopback =484;
13304: waveform_sig_loopback =1191;
13305: waveform_sig_loopback =2053;
13306: waveform_sig_loopback =1326;
13307: waveform_sig_loopback =1931;
13308: waveform_sig_loopback =186;
13309: waveform_sig_loopback =2271;
13310: waveform_sig_loopback =1496;
13311: waveform_sig_loopback =515;
13312: waveform_sig_loopback =1713;
13313: waveform_sig_loopback =998;
13314: waveform_sig_loopback =1252;
13315: waveform_sig_loopback =456;
13316: waveform_sig_loopback =2210;
13317: waveform_sig_loopback =178;
13318: waveform_sig_loopback =630;
13319: waveform_sig_loopback =1759;
13320: waveform_sig_loopback =638;
13321: waveform_sig_loopback =104;
13322: waveform_sig_loopback =1379;
13323: waveform_sig_loopback =1389;
13324: waveform_sig_loopback =-921;
13325: waveform_sig_loopback =1341;
13326: waveform_sig_loopback =1594;
13327: waveform_sig_loopback =-855;
13328: waveform_sig_loopback =322;
13329: waveform_sig_loopback =1531;
13330: waveform_sig_loopback =443;
13331: waveform_sig_loopback =-1025;
13332: waveform_sig_loopback =919;
13333: waveform_sig_loopback =1462;
13334: waveform_sig_loopback =-1364;
13335: waveform_sig_loopback =2242;
13336: waveform_sig_loopback =-2355;
13337: waveform_sig_loopback =-889;
13338: waveform_sig_loopback =3068;
13339: waveform_sig_loopback =-984;
13340: waveform_sig_loopback =-931;
13341: waveform_sig_loopback =-650;
13342: waveform_sig_loopback =461;
13343: waveform_sig_loopback =1009;
13344: waveform_sig_loopback =-1491;
13345: waveform_sig_loopback =-509;
13346: waveform_sig_loopback =320;
13347: waveform_sig_loopback =-962;
13348: waveform_sig_loopback =115;
13349: waveform_sig_loopback =-1353;
13350: waveform_sig_loopback =138;
13351: waveform_sig_loopback =-470;
13352: waveform_sig_loopback =-1319;
13353: waveform_sig_loopback =-201;
13354: waveform_sig_loopback =-874;
13355: waveform_sig_loopback =-817;
13356: waveform_sig_loopback =-1368;
13357: waveform_sig_loopback =368;
13358: waveform_sig_loopback =-1770;
13359: waveform_sig_loopback =-1506;
13360: waveform_sig_loopback =195;
13361: waveform_sig_loopback =-1468;
13362: waveform_sig_loopback =-1907;
13363: waveform_sig_loopback =-137;
13364: waveform_sig_loopback =-1113;
13365: waveform_sig_loopback =-2330;
13366: waveform_sig_loopback =-713;
13367: waveform_sig_loopback =-624;
13368: waveform_sig_loopback =-2239;
13369: waveform_sig_loopback =-1998;
13370: waveform_sig_loopback =-81;
13371: waveform_sig_loopback =-1524;
13372: waveform_sig_loopback =-3240;
13373: waveform_sig_loopback =-375;
13374: waveform_sig_loopback =-964;
13375: waveform_sig_loopback =-3077;
13376: waveform_sig_loopback =636;
13377: waveform_sig_loopback =-4834;
13378: waveform_sig_loopback =-2189;
13379: waveform_sig_loopback =1015;
13380: waveform_sig_loopback =-2834;
13381: waveform_sig_loopback =-2674;
13382: waveform_sig_loopback =-2805;
13383: waveform_sig_loopback =-1199;
13384: waveform_sig_loopback =-651;
13385: waveform_sig_loopback =-3697;
13386: waveform_sig_loopback =-2443;
13387: waveform_sig_loopback =-1460;
13388: waveform_sig_loopback =-2734;
13389: waveform_sig_loopback =-1803;
13390: waveform_sig_loopback =-3401;
13391: waveform_sig_loopback =-1641;
13392: waveform_sig_loopback =-2211;
13393: waveform_sig_loopback =-3215;
13394: waveform_sig_loopback =-2272;
13395: waveform_sig_loopback =-2403;
13396: waveform_sig_loopback =-2827;
13397: waveform_sig_loopback =-3231;
13398: waveform_sig_loopback =-1269;
13399: waveform_sig_loopback =-4072;
13400: waveform_sig_loopback =-2751;
13401: waveform_sig_loopback =-1877;
13402: waveform_sig_loopback =-3569;
13403: waveform_sig_loopback =-3224;
13404: waveform_sig_loopback =-2317;
13405: waveform_sig_loopback =-2773;
13406: waveform_sig_loopback =-4135;
13407: waveform_sig_loopback =-2649;
13408: waveform_sig_loopback =-2127;
13409: waveform_sig_loopback =-4327;
13410: waveform_sig_loopback =-3763;
13411: waveform_sig_loopback =-1654;
13412: waveform_sig_loopback =-3600;
13413: waveform_sig_loopback =-4907;
13414: waveform_sig_loopback =-1976;
13415: waveform_sig_loopback =-3096;
13416: waveform_sig_loopback =-4522;
13417: waveform_sig_loopback =-1239;
13418: waveform_sig_loopback =-6837;
13419: waveform_sig_loopback =-3470;
13420: waveform_sig_loopback =-968;
13421: waveform_sig_loopback =-4681;
13422: waveform_sig_loopback =-4243;
13423: waveform_sig_loopback =-4766;
13424: waveform_sig_loopback =-2673;
13425: waveform_sig_loopback =-2390;
13426: waveform_sig_loopback =-5617;
13427: waveform_sig_loopback =-3767;
13428: waveform_sig_loopback =-3380;
13429: waveform_sig_loopback =-4464;
13430: waveform_sig_loopback =-3225;
13431: waveform_sig_loopback =-5350;
13432: waveform_sig_loopback =-3162;
13433: waveform_sig_loopback =-3835;
13434: waveform_sig_loopback =-5051;
13435: waveform_sig_loopback =-3723;
13436: waveform_sig_loopback =-4097;
13437: waveform_sig_loopback =-4671;
13438: waveform_sig_loopback =-4507;
13439: waveform_sig_loopback =-3187;
13440: waveform_sig_loopback =-5716;
13441: waveform_sig_loopback =-4073;
13442: waveform_sig_loopback =-3916;
13443: waveform_sig_loopback =-4907;
13444: waveform_sig_loopback =-4897;
13445: waveform_sig_loopback =-4068;
13446: waveform_sig_loopback =-4096;
13447: waveform_sig_loopback =-6009;
13448: waveform_sig_loopback =-4032;
13449: waveform_sig_loopback =-3654;
13450: waveform_sig_loopback =-6193;
13451: waveform_sig_loopback =-5009;
13452: waveform_sig_loopback =-3244;
13453: waveform_sig_loopback =-5367;
13454: waveform_sig_loopback =-6263;
13455: waveform_sig_loopback =-3466;
13456: waveform_sig_loopback =-4864;
13457: waveform_sig_loopback =-5734;
13458: waveform_sig_loopback =-2996;
13459: waveform_sig_loopback =-8491;
13460: waveform_sig_loopback =-4470;
13461: waveform_sig_loopback =-2928;
13462: waveform_sig_loopback =-5951;
13463: waveform_sig_loopback =-5790;
13464: waveform_sig_loopback =-6325;
13465: waveform_sig_loopback =-3736;
13466: waveform_sig_loopback =-4270;
13467: waveform_sig_loopback =-7087;
13468: waveform_sig_loopback =-4913;
13469: waveform_sig_loopback =-5155;
13470: waveform_sig_loopback =-5558;
13471: waveform_sig_loopback =-4813;
13472: waveform_sig_loopback =-6887;
13473: waveform_sig_loopback =-4168;
13474: waveform_sig_loopback =-5591;
13475: waveform_sig_loopback =-6335;
13476: waveform_sig_loopback =-4937;
13477: waveform_sig_loopback =-5706;
13478: waveform_sig_loopback =-5885;
13479: waveform_sig_loopback =-5819;
13480: waveform_sig_loopback =-4689;
13481: waveform_sig_loopback =-6887;
13482: waveform_sig_loopback =-5460;
13483: waveform_sig_loopback =-5340;
13484: waveform_sig_loopback =-6045;
13485: waveform_sig_loopback =-6436;
13486: waveform_sig_loopback =-5173;
13487: waveform_sig_loopback =-5400;
13488: waveform_sig_loopback =-7566;
13489: waveform_sig_loopback =-4917;
13490: waveform_sig_loopback =-5103;
13491: waveform_sig_loopback =-7642;
13492: waveform_sig_loopback =-5836;
13493: waveform_sig_loopback =-4763;
13494: waveform_sig_loopback =-6597;
13495: waveform_sig_loopback =-7323;
13496: waveform_sig_loopback =-4863;
13497: waveform_sig_loopback =-5925;
13498: waveform_sig_loopback =-6913;
13499: waveform_sig_loopback =-4422;
13500: waveform_sig_loopback =-9489;
13501: waveform_sig_loopback =-5587;
13502: waveform_sig_loopback =-4168;
13503: waveform_sig_loopback =-6975;
13504: waveform_sig_loopback =-7223;
13505: waveform_sig_loopback =-7174;
13506: waveform_sig_loopback =-4806;
13507: waveform_sig_loopback =-5642;
13508: waveform_sig_loopback =-7938;
13509: waveform_sig_loopback =-6057;
13510: waveform_sig_loopback =-6331;
13511: waveform_sig_loopback =-6358;
13512: waveform_sig_loopback =-6181;
13513: waveform_sig_loopback =-7774;
13514: waveform_sig_loopback =-5074;
13515: waveform_sig_loopback =-6979;
13516: waveform_sig_loopback =-7026;
13517: waveform_sig_loopback =-6059;
13518: waveform_sig_loopback =-6837;
13519: waveform_sig_loopback =-6622;
13520: waveform_sig_loopback =-6970;
13521: waveform_sig_loopback =-5658;
13522: waveform_sig_loopback =-7695;
13523: waveform_sig_loopback =-6638;
13524: waveform_sig_loopback =-6008;
13525: waveform_sig_loopback =-7059;
13526: waveform_sig_loopback =-7463;
13527: waveform_sig_loopback =-5690;
13528: waveform_sig_loopback =-6704;
13529: waveform_sig_loopback =-8226;
13530: waveform_sig_loopback =-5600;
13531: waveform_sig_loopback =-6332;
13532: waveform_sig_loopback =-8195;
13533: waveform_sig_loopback =-6716;
13534: waveform_sig_loopback =-5658;
13535: waveform_sig_loopback =-7290;
13536: waveform_sig_loopback =-8215;
13537: waveform_sig_loopback =-5516;
13538: waveform_sig_loopback =-6710;
13539: waveform_sig_loopback =-7654;
13540: waveform_sig_loopback =-5186;
13541: waveform_sig_loopback =-10210;
13542: waveform_sig_loopback =-6245;
13543: waveform_sig_loopback =-4827;
13544: waveform_sig_loopback =-7773;
13545: waveform_sig_loopback =-8058;
13546: waveform_sig_loopback =-7486;
13547: waveform_sig_loopback =-5736;
13548: waveform_sig_loopback =-6271;
13549: waveform_sig_loopback =-8459;
13550: waveform_sig_loopback =-6945;
13551: waveform_sig_loopback =-6680;
13552: waveform_sig_loopback =-7121;
13553: waveform_sig_loopback =-6926;
13554: waveform_sig_loopback =-8000;
13555: waveform_sig_loopback =-5928;
13556: waveform_sig_loopback =-7515;
13557: waveform_sig_loopback =-7434;
13558: waveform_sig_loopback =-6832;
13559: waveform_sig_loopback =-7132;
13560: waveform_sig_loopback =-7268;
13561: waveform_sig_loopback =-7481;
13562: waveform_sig_loopback =-5956;
13563: waveform_sig_loopback =-8405;
13564: waveform_sig_loopback =-7026;
13565: waveform_sig_loopback =-6320;
13566: waveform_sig_loopback =-7802;
13567: waveform_sig_loopback =-7660;
13568: waveform_sig_loopback =-6099;
13569: waveform_sig_loopback =-7437;
13570: waveform_sig_loopback =-8261;
13571: waveform_sig_loopback =-6103;
13572: waveform_sig_loopback =-6841;
13573: waveform_sig_loopback =-8408;
13574: waveform_sig_loopback =-7176;
13575: waveform_sig_loopback =-5903;
13576: waveform_sig_loopback =-7729;
13577: waveform_sig_loopback =-8642;
13578: waveform_sig_loopback =-5557;
13579: waveform_sig_loopback =-7269;
13580: waveform_sig_loopback =-7913;
13581: waveform_sig_loopback =-5323;
13582: waveform_sig_loopback =-10767;
13583: waveform_sig_loopback =-6248;
13584: waveform_sig_loopback =-4988;
13585: waveform_sig_loopback =-8335;
13586: waveform_sig_loopback =-8071;
13587: waveform_sig_loopback =-7654;
13588: waveform_sig_loopback =-6095;
13589: waveform_sig_loopback =-6205;
13590: waveform_sig_loopback =-8959;
13591: waveform_sig_loopback =-6935;
13592: waveform_sig_loopback =-6709;
13593: waveform_sig_loopback =-7574;
13594: waveform_sig_loopback =-6811;
13595: waveform_sig_loopback =-8235;
13596: waveform_sig_loopback =-6110;
13597: waveform_sig_loopback =-7420;
13598: waveform_sig_loopback =-7663;
13599: waveform_sig_loopback =-6854;
13600: waveform_sig_loopback =-7093;
13601: waveform_sig_loopback =-7524;
13602: waveform_sig_loopback =-7347;
13603: waveform_sig_loopback =-6016;
13604: waveform_sig_loopback =-8580;
13605: waveform_sig_loopback =-6782;
13606: waveform_sig_loopback =-6408;
13607: waveform_sig_loopback =-7950;
13608: waveform_sig_loopback =-7338;
13609: waveform_sig_loopback =-6209;
13610: waveform_sig_loopback =-7467;
13611: waveform_sig_loopback =-7947;
13612: waveform_sig_loopback =-6254;
13613: waveform_sig_loopback =-6583;
13614: waveform_sig_loopback =-8365;
13615: waveform_sig_loopback =-7164;
13616: waveform_sig_loopback =-5461;
13617: waveform_sig_loopback =-7891;
13618: waveform_sig_loopback =-8388;
13619: waveform_sig_loopback =-5101;
13620: waveform_sig_loopback =-7527;
13621: waveform_sig_loopback =-7298;
13622: waveform_sig_loopback =-5325;
13623: waveform_sig_loopback =-10801;
13624: waveform_sig_loopback =-5414;
13625: waveform_sig_loopback =-5201;
13626: waveform_sig_loopback =-8046;
13627: waveform_sig_loopback =-7592;
13628: waveform_sig_loopback =-7667;
13629: waveform_sig_loopback =-5468;
13630: waveform_sig_loopback =-6091;
13631: waveform_sig_loopback =-8804;
13632: waveform_sig_loopback =-6197;
13633: waveform_sig_loopback =-6667;
13634: waveform_sig_loopback =-7072;
13635: waveform_sig_loopback =-6460;
13636: waveform_sig_loopback =-8002;
13637: waveform_sig_loopback =-5434;
13638: waveform_sig_loopback =-7224;
13639: waveform_sig_loopback =-7243;
13640: waveform_sig_loopback =-6423;
13641: waveform_sig_loopback =-6562;
13642: waveform_sig_loopback =-7306;
13643: waveform_sig_loopback =-6637;
13644: waveform_sig_loopback =-5642;
13645: waveform_sig_loopback =-8287;
13646: waveform_sig_loopback =-5839;
13647: waveform_sig_loopback =-6321;
13648: waveform_sig_loopback =-7209;
13649: waveform_sig_loopback =-6675;
13650: waveform_sig_loopback =-5994;
13651: waveform_sig_loopback =-6502;
13652: waveform_sig_loopback =-7707;
13653: waveform_sig_loopback =-5535;
13654: waveform_sig_loopback =-5793;
13655: waveform_sig_loopback =-8206;
13656: waveform_sig_loopback =-6055;
13657: waveform_sig_loopback =-5010;
13658: waveform_sig_loopback =-7447;
13659: waveform_sig_loopback =-7308;
13660: waveform_sig_loopback =-4723;
13661: waveform_sig_loopback =-6878;
13662: waveform_sig_loopback =-6335;
13663: waveform_sig_loopback =-4963;
13664: waveform_sig_loopback =-9908;
13665: waveform_sig_loopback =-4568;
13666: waveform_sig_loopback =-4685;
13667: waveform_sig_loopback =-7115;
13668: waveform_sig_loopback =-6951;
13669: waveform_sig_loopback =-6905;
13670: waveform_sig_loopback =-4451;
13671: waveform_sig_loopback =-5502;
13672: waveform_sig_loopback =-8018;
13673: waveform_sig_loopback =-5197;
13674: waveform_sig_loopback =-6183;
13675: waveform_sig_loopback =-5933;
13676: waveform_sig_loopback =-5666;
13677: waveform_sig_loopback =-7295;
13678: waveform_sig_loopback =-4343;
13679: waveform_sig_loopback =-6522;
13680: waveform_sig_loopback =-6356;
13681: waveform_sig_loopback =-5248;
13682: waveform_sig_loopback =-6016;
13683: waveform_sig_loopback =-6195;
13684: waveform_sig_loopback =-5515;
13685: waveform_sig_loopback =-5236;
13686: waveform_sig_loopback =-6842;
13687: waveform_sig_loopback =-5194;
13688: waveform_sig_loopback =-5364;
13689: waveform_sig_loopback =-6173;
13690: waveform_sig_loopback =-6092;
13691: waveform_sig_loopback =-4463;
13692: waveform_sig_loopback =-5758;
13693: waveform_sig_loopback =-6964;
13694: waveform_sig_loopback =-4231;
13695: waveform_sig_loopback =-4926;
13696: waveform_sig_loopback =-7099;
13697: waveform_sig_loopback =-4961;
13698: waveform_sig_loopback =-4193;
13699: waveform_sig_loopback =-6170;
13700: waveform_sig_loopback =-6181;
13701: waveform_sig_loopback =-3800;
13702: waveform_sig_loopback =-5749;
13703: waveform_sig_loopback =-5031;
13704: waveform_sig_loopback =-4130;
13705: waveform_sig_loopback =-8763;
13706: waveform_sig_loopback =-3204;
13707: waveform_sig_loopback =-3703;
13708: waveform_sig_loopback =-5897;
13709: waveform_sig_loopback =-6029;
13710: waveform_sig_loopback =-5555;
13711: waveform_sig_loopback =-3048;
13712: waveform_sig_loopback =-4764;
13713: waveform_sig_loopback =-6553;
13714: waveform_sig_loopback =-3990;
13715: waveform_sig_loopback =-5158;
13716: waveform_sig_loopback =-4377;
13717: waveform_sig_loopback =-4932;
13718: waveform_sig_loopback =-5696;
13719: waveform_sig_loopback =-3051;
13720: waveform_sig_loopback =-5714;
13721: waveform_sig_loopback =-4605;
13722: waveform_sig_loopback =-4205;
13723: waveform_sig_loopback =-4819;
13724: waveform_sig_loopback =-4642;
13725: waveform_sig_loopback =-4539;
13726: waveform_sig_loopback =-3647;
13727: waveform_sig_loopback =-5558;
13728: waveform_sig_loopback =-4005;
13729: waveform_sig_loopback =-3704;
13730: waveform_sig_loopback =-4990;
13731: waveform_sig_loopback =-4548;
13732: waveform_sig_loopback =-3117;
13733: waveform_sig_loopback =-4669;
13734: waveform_sig_loopback =-5092;
13735: waveform_sig_loopback =-2834;
13736: waveform_sig_loopback =-3873;
13737: waveform_sig_loopback =-5597;
13738: waveform_sig_loopback =-3249;
13739: waveform_sig_loopback =-2917;
13740: waveform_sig_loopback =-4965;
13741: waveform_sig_loopback =-4555;
13742: waveform_sig_loopback =-2383;
13743: waveform_sig_loopback =-4213;
13744: waveform_sig_loopback =-3614;
13745: waveform_sig_loopback =-2908;
13746: waveform_sig_loopback =-6875;
13747: waveform_sig_loopback =-1933;
13748: waveform_sig_loopback =-2117;
13749: waveform_sig_loopback =-4354;
13750: waveform_sig_loopback =-4756;
13751: waveform_sig_loopback =-3465;
13752: waveform_sig_loopback =-2011;
13753: waveform_sig_loopback =-3164;
13754: waveform_sig_loopback =-4725;
13755: waveform_sig_loopback =-2888;
13756: waveform_sig_loopback =-3200;
13757: waveform_sig_loopback =-2926;
13758: waveform_sig_loopback =-3466;
13759: waveform_sig_loopback =-3762;
13760: waveform_sig_loopback =-1886;
13761: waveform_sig_loopback =-3869;
13762: waveform_sig_loopback =-2934;
13763: waveform_sig_loopback =-2910;
13764: waveform_sig_loopback =-2782;
13765: waveform_sig_loopback =-3327;
13766: waveform_sig_loopback =-2662;
13767: waveform_sig_loopback =-2035;
13768: waveform_sig_loopback =-4097;
13769: waveform_sig_loopback =-2097;
13770: waveform_sig_loopback =-2175;
13771: waveform_sig_loopback =-3262;
13772: waveform_sig_loopback =-2941;
13773: waveform_sig_loopback =-1303;
13774: waveform_sig_loopback =-3170;
13775: waveform_sig_loopback =-3349;
13776: waveform_sig_loopback =-1010;
13777: waveform_sig_loopback =-2547;
13778: waveform_sig_loopback =-3504;
13779: waveform_sig_loopback =-1735;
13780: waveform_sig_loopback =-1267;
13781: waveform_sig_loopback =-2981;
13782: waveform_sig_loopback =-3213;
13783: waveform_sig_loopback =-229;
13784: waveform_sig_loopback =-2741;
13785: waveform_sig_loopback =-1944;
13786: waveform_sig_loopback =-865;
13787: waveform_sig_loopback =-5560;
13788: waveform_sig_loopback =232;
13789: waveform_sig_loopback =-350;
13790: waveform_sig_loopback =-3093;
13791: waveform_sig_loopback =-2482;
13792: waveform_sig_loopback =-1912;
13793: waveform_sig_loopback =-288;
13794: waveform_sig_loopback =-1108;
13795: waveform_sig_loopback =-3307;
13796: waveform_sig_loopback =-733;
13797: waveform_sig_loopback =-1476;
13798: waveform_sig_loopback =-1366;
13799: waveform_sig_loopback =-1413;
13800: waveform_sig_loopback =-2047;
13801: waveform_sig_loopback =-109;
13802: waveform_sig_loopback =-1941;
13803: waveform_sig_loopback =-1288;
13804: waveform_sig_loopback =-979;
13805: waveform_sig_loopback =-983;
13806: waveform_sig_loopback =-1626;
13807: waveform_sig_loopback =-709;
13808: waveform_sig_loopback =-248;
13809: waveform_sig_loopback =-2314;
13810: waveform_sig_loopback =-181;
13811: waveform_sig_loopback =-316;
13812: waveform_sig_loopback =-1702;
13813: waveform_sig_loopback =-735;
13814: waveform_sig_loopback =358;
13815: waveform_sig_loopback =-1528;
13816: waveform_sig_loopback =-1056;
13817: waveform_sig_loopback =485;
13818: waveform_sig_loopback =-503;
13819: waveform_sig_loopback =-1655;
13820: waveform_sig_loopback =-77;
13821: waveform_sig_loopback =999;
13822: waveform_sig_loopback =-1556;
13823: waveform_sig_loopback =-1167;
13824: waveform_sig_loopback =1941;
13825: waveform_sig_loopback =-1514;
13826: waveform_sig_loopback =572;
13827: waveform_sig_loopback =625;
13828: waveform_sig_loopback =-3790;
13829: waveform_sig_loopback =2737;
13830: waveform_sig_loopback =844;
13831: waveform_sig_loopback =-964;
13832: waveform_sig_loopback =-544;
13833: waveform_sig_loopback =-304;
13834: waveform_sig_loopback =1998;
13835: waveform_sig_loopback =359;
13836: waveform_sig_loopback =-1381;
13837: waveform_sig_loopback =1347;
13838: waveform_sig_loopback =171;
13839: waveform_sig_loopback =712;
13840: waveform_sig_loopback =339;
13841: waveform_sig_loopback =-142;
13842: waveform_sig_loopback =1839;
13843: waveform_sig_loopback =-78;
13844: waveform_sig_loopback =609;
13845: waveform_sig_loopback =836;
13846: waveform_sig_loopback =1106;
13847: waveform_sig_loopback =-61;
13848: waveform_sig_loopback =1485;
13849: waveform_sig_loopback =1445;
13850: waveform_sig_loopback =-584;
13851: waveform_sig_loopback =2227;
13852: waveform_sig_loopback =929;
13853: waveform_sig_loopback =532;
13854: waveform_sig_loopback =1259;
13855: waveform_sig_loopback =1866;
13856: waveform_sig_loopback =826;
13857: waveform_sig_loopback =417;
13858: waveform_sig_loopback =2597;
13859: waveform_sig_loopback =1412;
13860: waveform_sig_loopback =-119;
13861: waveform_sig_loopback =2312;
13862: waveform_sig_loopback =2593;
13863: waveform_sig_loopback =139;
13864: waveform_sig_loopback =1091;
13865: waveform_sig_loopback =3527;
13866: waveform_sig_loopback =340;
13867: waveform_sig_loopback =2698;
13868: waveform_sig_loopback =1963;
13869: waveform_sig_loopback =-1622;
13870: waveform_sig_loopback =4645;
13871: waveform_sig_loopback =2433;
13872: waveform_sig_loopback =1134;
13873: waveform_sig_loopback =1130;
13874: waveform_sig_loopback =1644;
13875: waveform_sig_loopback =4074;
13876: waveform_sig_loopback =1949;
13877: waveform_sig_loopback =604;
13878: waveform_sig_loopback =3305;
13879: waveform_sig_loopback =1812;
13880: waveform_sig_loopback =2862;
13881: waveform_sig_loopback =2065;
13882: waveform_sig_loopback =1642;
13883: waveform_sig_loopback =3924;
13884: waveform_sig_loopback =1563;
13885: waveform_sig_loopback =2487;
13886: waveform_sig_loopback =2871;
13887: waveform_sig_loopback =2684;
13888: waveform_sig_loopback =1933;
13889: waveform_sig_loopback =3471;
13890: waveform_sig_loopback =2812;
13891: waveform_sig_loopback =1704;
13892: waveform_sig_loopback =3798;
13893: waveform_sig_loopback =2667;
13894: waveform_sig_loopback =2610;
13895: waveform_sig_loopback =2624;
13896: waveform_sig_loopback =3991;
13897: waveform_sig_loopback =2419;
13898: waveform_sig_loopback =2099;
13899: waveform_sig_loopback =4674;
13900: waveform_sig_loopback =2821;
13901: waveform_sig_loopback =1754;
13902: waveform_sig_loopback =4209;
13903: waveform_sig_loopback =4136;
13904: waveform_sig_loopback =1967;
13905: waveform_sig_loopback =3037;
13906: waveform_sig_loopback =5121;
13907: waveform_sig_loopback =2168;
13908: waveform_sig_loopback =4647;
13909: waveform_sig_loopback =3361;
13910: waveform_sig_loopback =540;
13911: waveform_sig_loopback =6356;
13912: waveform_sig_loopback =4084;
13913: waveform_sig_loopback =3066;
13914: waveform_sig_loopback =2587;
13915: waveform_sig_loopback =3756;
13916: waveform_sig_loopback =5725;
13917: waveform_sig_loopback =3375;
13918: waveform_sig_loopback =2642;
13919: waveform_sig_loopback =4919;
13920: waveform_sig_loopback =3445;
13921: waveform_sig_loopback =4722;
13922: waveform_sig_loopback =3473;
13923: waveform_sig_loopback =3530;
13924: waveform_sig_loopback =5638;
13925: waveform_sig_loopback =2909;
13926: waveform_sig_loopback =4434;
13927: waveform_sig_loopback =4407;
13928: waveform_sig_loopback =4125;
13929: waveform_sig_loopback =3830;
13930: waveform_sig_loopback =4850;
13931: waveform_sig_loopback =4509;
13932: waveform_sig_loopback =3446;
13933: waveform_sig_loopback =5079;
13934: waveform_sig_loopback =4654;
13935: waveform_sig_loopback =4024;
13936: waveform_sig_loopback =4221;
13937: waveform_sig_loopback =5820;
13938: waveform_sig_loopback =3638;
13939: waveform_sig_loopback =3967;
13940: waveform_sig_loopback =6297;
13941: waveform_sig_loopback =4146;
13942: waveform_sig_loopback =3553;
13943: waveform_sig_loopback =5829;
13944: waveform_sig_loopback =5569;
13945: waveform_sig_loopback =3616;
13946: waveform_sig_loopback =4581;
13947: waveform_sig_loopback =6633;
13948: waveform_sig_loopback =3808;
13949: waveform_sig_loopback =6107;
13950: waveform_sig_loopback =4716;
13951: waveform_sig_loopback =2251;
13952: waveform_sig_loopback =7743;
13953: waveform_sig_loopback =5634;
13954: waveform_sig_loopback =4363;
13955: waveform_sig_loopback =4017;
13956: waveform_sig_loopback =5515;
13957: waveform_sig_loopback =6858;
13958: waveform_sig_loopback =4879;
13959: waveform_sig_loopback =4187;
13960: waveform_sig_loopback =6109;
13961: waveform_sig_loopback =5041;
13962: waveform_sig_loopback =6017;
13963: waveform_sig_loopback =4709;
13964: waveform_sig_loopback =5260;
13965: waveform_sig_loopback =6726;
13966: waveform_sig_loopback =4353;
13967: waveform_sig_loopback =5991;
13968: waveform_sig_loopback =5538;
13969: waveform_sig_loopback =5702;
13970: waveform_sig_loopback =5168;
13971: waveform_sig_loopback =6151;
13972: waveform_sig_loopback =6003;
13973: waveform_sig_loopback =4653;
13974: waveform_sig_loopback =6466;
13975: waveform_sig_loopback =6129;
13976: waveform_sig_loopback =4940;
13977: waveform_sig_loopback =5929;
13978: waveform_sig_loopback =7070;
13979: waveform_sig_loopback =4628;
13980: waveform_sig_loopback =5674;
13981: waveform_sig_loopback =7292;
13982: waveform_sig_loopback =5393;
13983: waveform_sig_loopback =5057;
13984: waveform_sig_loopback =6816;
13985: waveform_sig_loopback =6908;
13986: waveform_sig_loopback =4746;
13987: waveform_sig_loopback =5804;
13988: waveform_sig_loopback =7928;
13989: waveform_sig_loopback =4734;
13990: waveform_sig_loopback =7428;
13991: waveform_sig_loopback =5826;
13992: waveform_sig_loopback =3340;
13993: waveform_sig_loopback =9059;
13994: waveform_sig_loopback =6727;
13995: waveform_sig_loopback =5229;
13996: waveform_sig_loopback =5354;
13997: waveform_sig_loopback =6632;
13998: waveform_sig_loopback =7840;
13999: waveform_sig_loopback =6069;
14000: waveform_sig_loopback =5161;
14001: waveform_sig_loopback =7241;
14002: waveform_sig_loopback =6272;
14003: waveform_sig_loopback =6800;
14004: waveform_sig_loopback =5875;
14005: waveform_sig_loopback =6465;
14006: waveform_sig_loopback =7417;
14007: waveform_sig_loopback =5693;
14008: waveform_sig_loopback =6839;
14009: waveform_sig_loopback =6487;
14010: waveform_sig_loopback =6998;
14011: waveform_sig_loopback =5748;
14012: waveform_sig_loopback =7488;
14013: waveform_sig_loopback =6877;
14014: waveform_sig_loopback =5388;
14015: waveform_sig_loopback =7855;
14016: waveform_sig_loopback =6667;
14017: waveform_sig_loopback =5971;
14018: waveform_sig_loopback =7063;
14019: waveform_sig_loopback =7582;
14020: waveform_sig_loopback =5745;
14021: waveform_sig_loopback =6556;
14022: waveform_sig_loopback =8068;
14023: waveform_sig_loopback =6273;
14024: waveform_sig_loopback =5808;
14025: waveform_sig_loopback =7797;
14026: waveform_sig_loopback =7660;
14027: waveform_sig_loopback =5445;
14028: waveform_sig_loopback =6617;
14029: waveform_sig_loopback =8859;
14030: waveform_sig_loopback =5274;
14031: waveform_sig_loopback =8397;
14032: waveform_sig_loopback =6357;
14033: waveform_sig_loopback =4073;
14034: waveform_sig_loopback =10142;
14035: waveform_sig_loopback =7127;
14036: waveform_sig_loopback =5887;
14037: waveform_sig_loopback =6334;
14038: waveform_sig_loopback =7079;
14039: waveform_sig_loopback =8708;
14040: waveform_sig_loopback =6580;
14041: waveform_sig_loopback =5481;
14042: waveform_sig_loopback =8403;
14043: waveform_sig_loopback =6632;
14044: waveform_sig_loopback =7397;
14045: waveform_sig_loopback =6464;
14046: waveform_sig_loopback =6971;
14047: waveform_sig_loopback =8319;
14048: waveform_sig_loopback =6065;
14049: waveform_sig_loopback =7179;
14050: waveform_sig_loopback =7357;
14051: waveform_sig_loopback =7387;
14052: waveform_sig_loopback =6181;
14053: waveform_sig_loopback =8141;
14054: waveform_sig_loopback =7159;
14055: waveform_sig_loopback =6044;
14056: waveform_sig_loopback =8306;
14057: waveform_sig_loopback =6914;
14058: waveform_sig_loopback =6597;
14059: waveform_sig_loopback =7499;
14060: waveform_sig_loopback =7777;
14061: waveform_sig_loopback =6286;
14062: waveform_sig_loopback =6970;
14063: waveform_sig_loopback =8421;
14064: waveform_sig_loopback =6679;
14065: waveform_sig_loopback =5987;
14066: waveform_sig_loopback =8352;
14067: waveform_sig_loopback =7980;
14068: waveform_sig_loopback =5476;
14069: waveform_sig_loopback =7358;
14070: waveform_sig_loopback =8956;
14071: waveform_sig_loopback =5443;
14072: waveform_sig_loopback =9052;
14073: waveform_sig_loopback =6107;
14074: waveform_sig_loopback =4679;
14075: waveform_sig_loopback =10535;
14076: waveform_sig_loopback =6917;
14077: waveform_sig_loopback =6517;
14078: waveform_sig_loopback =6389;
14079: waveform_sig_loopback =7172;
14080: waveform_sig_loopback =9230;
14081: waveform_sig_loopback =6363;
14082: waveform_sig_loopback =6070;
14083: waveform_sig_loopback =8439;
14084: waveform_sig_loopback =6401;
14085: waveform_sig_loopback =8069;
14086: waveform_sig_loopback =6429;
14087: waveform_sig_loopback =7007;
14088: waveform_sig_loopback =8452;
14089: waveform_sig_loopback =5974;
14090: waveform_sig_loopback =7579;
14091: waveform_sig_loopback =7294;
14092: waveform_sig_loopback =7157;
14093: waveform_sig_loopback =6514;
14094: waveform_sig_loopback =8215;
14095: waveform_sig_loopback =6858;
14096: waveform_sig_loopback =6238;
14097: waveform_sig_loopback =8301;
14098: waveform_sig_loopback =6809;
14099: waveform_sig_loopback =6630;
14100: waveform_sig_loopback =7385;
14101: waveform_sig_loopback =7766;
14102: waveform_sig_loopback =6349;
14103: waveform_sig_loopback =6640;
14104: waveform_sig_loopback =8535;
14105: waveform_sig_loopback =6555;
14106: waveform_sig_loopback =5646;
14107: waveform_sig_loopback =8695;
14108: waveform_sig_loopback =7371;
14109: waveform_sig_loopback =5450;
14110: waveform_sig_loopback =7540;
14111: waveform_sig_loopback =8204;
14112: waveform_sig_loopback =5754;
14113: waveform_sig_loopback =8736;
14114: waveform_sig_loopback =5529;
14115: waveform_sig_loopback =5001;
14116: waveform_sig_loopback =9884;
14117: waveform_sig_loopback =6886;
14118: waveform_sig_loopback =6229;
14119: waveform_sig_loopback =5782;
14120: waveform_sig_loopback =7351;
14121: waveform_sig_loopback =8748;
14122: waveform_sig_loopback =5924;
14123: waveform_sig_loopback =5982;
14124: waveform_sig_loopback =7924;
14125: waveform_sig_loopback =6158;
14126: waveform_sig_loopback =7790;
14127: waveform_sig_loopback =5809;
14128: waveform_sig_loopback =6887;
14129: waveform_sig_loopback =8012;
14130: waveform_sig_loopback =5447;
14131: waveform_sig_loopback =7335;
14132: waveform_sig_loopback =6801;
14133: waveform_sig_loopback =6576;
14134: waveform_sig_loopback =6291;
14135: waveform_sig_loopback =7608;
14136: waveform_sig_loopback =6224;
14137: waveform_sig_loopback =6104;
14138: waveform_sig_loopback =7397;
14139: waveform_sig_loopback =6571;
14140: waveform_sig_loopback =6008;
14141: waveform_sig_loopback =6706;
14142: waveform_sig_loopback =7612;
14143: waveform_sig_loopback =5284;
14144: waveform_sig_loopback =6373;
14145: waveform_sig_loopback =8039;
14146: waveform_sig_loopback =5530;
14147: waveform_sig_loopback =5492;
14148: waveform_sig_loopback =7877;
14149: waveform_sig_loopback =6623;
14150: waveform_sig_loopback =5054;
14151: waveform_sig_loopback =6731;
14152: waveform_sig_loopback =7631;
14153: waveform_sig_loopback =5116;
14154: waveform_sig_loopback =8026;
14155: waveform_sig_loopback =4765;
14156: waveform_sig_loopback =4471;
14157: waveform_sig_loopback =9140;
14158: waveform_sig_loopback =6148;
14159: waveform_sig_loopback =5399;
14160: waveform_sig_loopback =5082;
14161: waveform_sig_loopback =6796;
14162: waveform_sig_loopback =7741;
14163: waveform_sig_loopback =5076;
14164: waveform_sig_loopback =5453;
14165: waveform_sig_loopback =6840;
14166: waveform_sig_loopback =5558;
14167: waveform_sig_loopback =6918;
14168: waveform_sig_loopback =4759;
14169: waveform_sig_loopback =6462;
14170: waveform_sig_loopback =6738;
14171: waveform_sig_loopback =4706;
14172: waveform_sig_loopback =6678;
14173: waveform_sig_loopback =5590;
14174: waveform_sig_loopback =5974;
14175: waveform_sig_loopback =5315;
14176: waveform_sig_loopback =6592;
14177: waveform_sig_loopback =5541;
14178: waveform_sig_loopback =4932;
14179: waveform_sig_loopback =6602;
14180: waveform_sig_loopback =5712;
14181: waveform_sig_loopback =4748;
14182: waveform_sig_loopback =6073;
14183: waveform_sig_loopback =6413;
14184: waveform_sig_loopback =4186;
14185: waveform_sig_loopback =5692;
14186: waveform_sig_loopback =6776;
14187: waveform_sig_loopback =4498;
14188: waveform_sig_loopback =4650;
14189: waveform_sig_loopback =6717;
14190: waveform_sig_loopback =5578;
14191: waveform_sig_loopback =4010;
14192: waveform_sig_loopback =5643;
14193: waveform_sig_loopback =6612;
14194: waveform_sig_loopback =3930;
14195: waveform_sig_loopback =6944;
14196: waveform_sig_loopback =3572;
14197: waveform_sig_loopback =3427;
14198: waveform_sig_loopback =8026;
14199: waveform_sig_loopback =5016;
14200: waveform_sig_loopback =4033;
14201: waveform_sig_loopback =4067;
14202: waveform_sig_loopback =5772;
14203: waveform_sig_loopback =6322;
14204: waveform_sig_loopback =4096;
14205: waveform_sig_loopback =4180;
14206: waveform_sig_loopback =5536;
14207: waveform_sig_loopback =4615;
14208: waveform_sig_loopback =5273;
14209: waveform_sig_loopback =3786;
14210: waveform_sig_loopback =5269;
14211: waveform_sig_loopback =5157;
14212: waveform_sig_loopback =3862;
14213: waveform_sig_loopback =5008;
14214: waveform_sig_loopback =4392;
14215: waveform_sig_loopback =4804;
14216: waveform_sig_loopback =3718;
14217: waveform_sig_loopback =5674;
14218: waveform_sig_loopback =3907;
14219: waveform_sig_loopback =3593;
14220: waveform_sig_loopback =5487;
14221: waveform_sig_loopback =4074;
14222: waveform_sig_loopback =3583;
14223: waveform_sig_loopback =4748;
14224: waveform_sig_loopback =4967;
14225: waveform_sig_loopback =2874;
14226: waveform_sig_loopback =4360;
14227: waveform_sig_loopback =5301;
14228: waveform_sig_loopback =2996;
14229: waveform_sig_loopback =3470;
14230: waveform_sig_loopback =5104;
14231: waveform_sig_loopback =4265;
14232: waveform_sig_loopback =2494;
14233: waveform_sig_loopback =4158;
14234: waveform_sig_loopback =5394;
14235: waveform_sig_loopback =2047;
14236: waveform_sig_loopback =5800;
14237: waveform_sig_loopback =1924;
14238: waveform_sig_loopback =1833;
14239: waveform_sig_loopback =6984;
14240: waveform_sig_loopback =3046;
14241: waveform_sig_loopback =2533;
14242: waveform_sig_loopback =2893;
14243: waveform_sig_loopback =3824;
14244: waveform_sig_loopback =5101;
14245: waveform_sig_loopback =2322;
14246: waveform_sig_loopback =2492;
14247: waveform_sig_loopback =4397;
14248: waveform_sig_loopback =2670;
14249: waveform_sig_loopback =3839;
14250: waveform_sig_loopback =2323;
14251: waveform_sig_loopback =3490;
14252: waveform_sig_loopback =3743;
14253: waveform_sig_loopback =2110;
14254: waveform_sig_loopback =3421;
14255: waveform_sig_loopback =2986;
14256: waveform_sig_loopback =2969;
14257: waveform_sig_loopback =2117;
14258: waveform_sig_loopback =4090;
14259: waveform_sig_loopback =2251;
14260: waveform_sig_loopback =2012;
14261: waveform_sig_loopback =3848;
14262: waveform_sig_loopback =2320;
14263: waveform_sig_loopback =1993;
14264: waveform_sig_loopback =3316;
14265: waveform_sig_loopback =2728;
14266: waveform_sig_loopback =1479;
14267: waveform_sig_loopback =2868;
14268: waveform_sig_loopback =3260;
14269: waveform_sig_loopback =1546;
14270: waveform_sig_loopback =1478;
14271: waveform_sig_loopback =3663;
14272: waveform_sig_loopback =2529;
14273: waveform_sig_loopback =279;
14274: waveform_sig_loopback =3085;
14275: waveform_sig_loopback =3219;
14276: waveform_sig_loopback =331;
14277: waveform_sig_loopback =4423;
14278: waveform_sig_loopback =-537;
14279: waveform_sig_loopback =746;
14280: waveform_sig_loopback =5106;
14281: waveform_sig_loopback =961;
14282: waveform_sig_loopback =1209;
14283: waveform_sig_loopback =884;
14284: waveform_sig_loopback =2195;
14285: waveform_sig_loopback =3404;
14286: waveform_sig_loopback =242;
14287: waveform_sig_loopback =1012;
14288: waveform_sig_loopback =2525;
14289: waveform_sig_loopback =746;
14290: waveform_sig_loopback =2247;
14291: waveform_sig_loopback =351;
14292: waveform_sig_loopback =1708;
14293: waveform_sig_loopback =1976;
14294: waveform_sig_loopback =301;
14295: waveform_sig_loopback =1545;
14296: waveform_sig_loopback =1259;
14297: waveform_sig_loopback =1023;
14298: waveform_sig_loopback =386;
14299: waveform_sig_loopback =2420;
14300: waveform_sig_loopback =-65;
14301: waveform_sig_loopback =631;
14302: waveform_sig_loopback =1982;
14303: waveform_sig_loopback =106;
14304: waveform_sig_loopback =603;
14305: waveform_sig_loopback =1148;
14306: waveform_sig_loopback =1041;
14307: waveform_sig_loopback =-240;
14308: waveform_sig_loopback =625;
14309: waveform_sig_loopback =1892;
14310: waveform_sig_loopback =-550;
14311: waveform_sig_loopback =-462;
14312: waveform_sig_loopback =2186;
14313: waveform_sig_loopback =188;
14314: waveform_sig_loopback =-1293;
14315: waveform_sig_loopback =1427;
14316: waveform_sig_loopback =824;
14317: waveform_sig_loopback =-1004;
14318: waveform_sig_loopback =2384;
14319: waveform_sig_loopback =-2749;
14320: waveform_sig_loopback =-512;
14321: waveform_sig_loopback =2769;
14322: waveform_sig_loopback =-775;
14323: waveform_sig_loopback =-660;
14324: waveform_sig_loopback =-1300;
14325: waveform_sig_loopback =748;
14326: waveform_sig_loopback =1338;
14327: waveform_sig_loopback =-1868;
14328: waveform_sig_loopback =-549;
14329: waveform_sig_loopback =416;
14330: waveform_sig_loopback =-1063;
14331: waveform_sig_loopback =473;
14332: waveform_sig_loopback =-1796;
14333: waveform_sig_loopback =74;
14334: waveform_sig_loopback =90;
14335: waveform_sig_loopback =-1838;
14336: waveform_sig_loopback =-93;
14337: waveform_sig_loopback =-588;
14338: waveform_sig_loopback =-1166;
14339: waveform_sig_loopback =-1027;
14340: waveform_sig_loopback =151;
14341: waveform_sig_loopback =-1870;
14342: waveform_sig_loopback =-873;
14343: waveform_sig_loopback =-506;
14344: waveform_sig_loopback =-1240;
14345: waveform_sig_loopback =-1535;
14346: waveform_sig_loopback =-798;
14347: waveform_sig_loopback =-436;
14348: waveform_sig_loopback =-2672;
14349: waveform_sig_loopback =-889;
14350: waveform_sig_loopback =45;
14351: waveform_sig_loopback =-2805;
14352: waveform_sig_loopback =-1882;
14353: waveform_sig_loopback =115;
14354: waveform_sig_loopback =-1759;
14355: waveform_sig_loopback =-2949;
14356: waveform_sig_loopback =-621;
14357: waveform_sig_loopback =-1005;
14358: waveform_sig_loopback =-2707;
14359: waveform_sig_loopback =318;
14360: waveform_sig_loopback =-4712;
14361: waveform_sig_loopback =-2036;
14362: waveform_sig_loopback =685;
14363: waveform_sig_loopback =-2559;
14364: waveform_sig_loopback =-2579;
14365: waveform_sig_loopback =-3273;
14366: waveform_sig_loopback =-682;
14367: waveform_sig_loopback =-875;
14368: waveform_sig_loopback =-3672;
14369: waveform_sig_loopback =-2074;
14370: waveform_sig_loopback =-1874;
14371: waveform_sig_loopback =-2519;
14372: waveform_sig_loopback =-1542;
14373: waveform_sig_loopback =-3785;
14374: waveform_sig_loopback =-1309;
14375: waveform_sig_loopback =-2190;
14376: waveform_sig_loopback =-3475;
14377: waveform_sig_loopback =-1760;
14378: waveform_sig_loopback =-2826;
14379: waveform_sig_loopback =-2674;
14380: waveform_sig_loopback =-2955;
14381: waveform_sig_loopback =-1833;
14382: waveform_sig_loopback =-3495;
14383: waveform_sig_loopback =-2853;
14384: waveform_sig_loopback =-2349;
14385: waveform_sig_loopback =-2899;
14386: waveform_sig_loopback =-3744;
14387: waveform_sig_loopback =-2331;
14388: waveform_sig_loopback =-2334;
14389: waveform_sig_loopback =-4747;
14390: waveform_sig_loopback =-2376;
14391: waveform_sig_loopback =-2219;
14392: waveform_sig_loopback =-4455;
14393: waveform_sig_loopback =-3344;
14394: waveform_sig_loopback =-2214;
14395: waveform_sig_loopback =-3562;
14396: waveform_sig_loopback =-4475;
14397: waveform_sig_loopback =-2475;
14398: waveform_sig_loopback =-2856;
14399: waveform_sig_loopback =-4608;
14400: waveform_sig_loopback =-1366;
14401: waveform_sig_loopback =-6344;
14402: waveform_sig_loopback =-3897;
14403: waveform_sig_loopback =-1129;
14404: waveform_sig_loopback =-4148;
14405: waveform_sig_loopback =-4575;
14406: waveform_sig_loopback =-4762;
14407: waveform_sig_loopback =-2437;
14408: waveform_sig_loopback =-2840;
14409: waveform_sig_loopback =-5161;
14410: waveform_sig_loopback =-3967;
14411: waveform_sig_loopback =-3655;
14412: waveform_sig_loopback =-3922;
14413: waveform_sig_loopback =-3669;
14414: waveform_sig_loopback =-5280;
14415: waveform_sig_loopback =-2919;
14416: waveform_sig_loopback =-4260;
14417: waveform_sig_loopback =-4755;
14418: waveform_sig_loopback =-3710;
14419: waveform_sig_loopback =-4535;
14420: waveform_sig_loopback =-4024;
14421: waveform_sig_loopback =-4944;
14422: waveform_sig_loopback =-3267;
14423: waveform_sig_loopback =-5132;
14424: waveform_sig_loopback =-4737;
14425: waveform_sig_loopback =-3564;
14426: waveform_sig_loopback =-4848;
14427: waveform_sig_loopback =-5292;
14428: waveform_sig_loopback =-3561;
14429: waveform_sig_loopback =-4409;
14430: waveform_sig_loopback =-6066;
14431: waveform_sig_loopback =-3704;
14432: waveform_sig_loopback =-4077;
14433: waveform_sig_loopback =-5974;
14434: waveform_sig_loopback =-4879;
14435: waveform_sig_loopback =-3658;
14436: waveform_sig_loopback =-4917;
14437: waveform_sig_loopback =-6384;
14438: waveform_sig_loopback =-3818;
14439: waveform_sig_loopback =-4230;
14440: waveform_sig_loopback =-6234;
14441: waveform_sig_loopback =-2917;
14442: waveform_sig_loopback =-8025;
14443: waveform_sig_loopback =-5205;
14444: waveform_sig_loopback =-2453;
14445: waveform_sig_loopback =-5912;
14446: waveform_sig_loopback =-6191;
14447: waveform_sig_loopback =-5795;
14448: waveform_sig_loopback =-4176;
14449: waveform_sig_loopback =-4298;
14450: waveform_sig_loopback =-6532;
14451: waveform_sig_loopback =-5563;
14452: waveform_sig_loopback =-4746;
14453: waveform_sig_loopback =-5584;
14454: waveform_sig_loopback =-5178;
14455: waveform_sig_loopback =-6309;
14456: waveform_sig_loopback =-4615;
14457: waveform_sig_loopback =-5569;
14458: waveform_sig_loopback =-5920;
14459: waveform_sig_loopback =-5372;
14460: waveform_sig_loopback =-5572;
14461: waveform_sig_loopback =-5608;
14462: waveform_sig_loopback =-6364;
14463: waveform_sig_loopback =-4252;
14464: waveform_sig_loopback =-6935;
14465: waveform_sig_loopback =-5897;
14466: waveform_sig_loopback =-4706;
14467: waveform_sig_loopback =-6573;
14468: waveform_sig_loopback =-6237;
14469: waveform_sig_loopback =-4988;
14470: waveform_sig_loopback =-5931;
14471: waveform_sig_loopback =-6940;
14472: waveform_sig_loopback =-5233;
14473: waveform_sig_loopback =-5245;
14474: waveform_sig_loopback =-7189;
14475: waveform_sig_loopback =-6304;
14476: waveform_sig_loopback =-4641;
14477: waveform_sig_loopback =-6379;
14478: waveform_sig_loopback =-7631;
14479: waveform_sig_loopback =-4762;
14480: waveform_sig_loopback =-5668;
14481: waveform_sig_loopback =-7345;
14482: waveform_sig_loopback =-4013;
14483: waveform_sig_loopback =-9445;
14484: waveform_sig_loopback =-6107;
14485: waveform_sig_loopback =-3506;
14486: waveform_sig_loopback =-7418;
14487: waveform_sig_loopback =-7102;
14488: waveform_sig_loopback =-6831;
14489: waveform_sig_loopback =-5559;
14490: waveform_sig_loopback =-4959;
14491: waveform_sig_loopback =-8086;
14492: waveform_sig_loopback =-6492;
14493: waveform_sig_loopback =-5585;
14494: waveform_sig_loopback =-7082;
14495: waveform_sig_loopback =-5776;
14496: waveform_sig_loopback =-7538;
14497: waveform_sig_loopback =-5767;
14498: waveform_sig_loopback =-6243;
14499: waveform_sig_loopback =-7323;
14500: waveform_sig_loopback =-6184;
14501: waveform_sig_loopback =-6405;
14502: waveform_sig_loopback =-7018;
14503: waveform_sig_loopback =-6832;
14504: waveform_sig_loopback =-5459;
14505: waveform_sig_loopback =-7970;
14506: waveform_sig_loopback =-6441;
14507: waveform_sig_loopback =-5983;
14508: waveform_sig_loopback =-7328;
14509: waveform_sig_loopback =-7088;
14510: waveform_sig_loopback =-5941;
14511: waveform_sig_loopback =-6803;
14512: waveform_sig_loopback =-7784;
14513: waveform_sig_loopback =-6125;
14514: waveform_sig_loopback =-6092;
14515: waveform_sig_loopback =-7959;
14516: waveform_sig_loopback =-7270;
14517: waveform_sig_loopback =-5200;
14518: waveform_sig_loopback =-7354;
14519: waveform_sig_loopback =-8469;
14520: waveform_sig_loopback =-5145;
14521: waveform_sig_loopback =-6998;
14522: waveform_sig_loopback =-7694;
14523: waveform_sig_loopback =-4783;
14524: waveform_sig_loopback =-10678;
14525: waveform_sig_loopback =-6046;
14526: waveform_sig_loopback =-4702;
14527: waveform_sig_loopback =-8166;
14528: waveform_sig_loopback =-7389;
14529: waveform_sig_loopback =-8032;
14530: waveform_sig_loopback =-5713;
14531: waveform_sig_loopback =-5743;
14532: waveform_sig_loopback =-9075;
14533: waveform_sig_loopback =-6470;
14534: waveform_sig_loopback =-6809;
14535: waveform_sig_loopback =-7456;
14536: waveform_sig_loopback =-6240;
14537: waveform_sig_loopback =-8576;
14538: waveform_sig_loopback =-5810;
14539: waveform_sig_loopback =-7177;
14540: waveform_sig_loopback =-7889;
14541: waveform_sig_loopback =-6499;
14542: waveform_sig_loopback =-7222;
14543: waveform_sig_loopback =-7387;
14544: waveform_sig_loopback =-7294;
14545: waveform_sig_loopback =-6098;
14546: waveform_sig_loopback =-8438;
14547: waveform_sig_loopback =-6795;
14548: waveform_sig_loopback =-6581;
14549: waveform_sig_loopback =-7767;
14550: waveform_sig_loopback =-7359;
14551: waveform_sig_loopback =-6594;
14552: waveform_sig_loopback =-6997;
14553: waveform_sig_loopback =-8307;
14554: waveform_sig_loopback =-6608;
14555: waveform_sig_loopback =-6140;
14556: waveform_sig_loopback =-8785;
14557: waveform_sig_loopback =-7266;
14558: waveform_sig_loopback =-5463;
14559: waveform_sig_loopback =-8240;
14560: waveform_sig_loopback =-8206;
14561: waveform_sig_loopback =-5683;
14562: waveform_sig_loopback =-7480;
14563: waveform_sig_loopback =-7429;
14564: waveform_sig_loopback =-5689;
14565: waveform_sig_loopback =-10640;
14566: waveform_sig_loopback =-6069;
14567: waveform_sig_loopback =-5447;
14568: waveform_sig_loopback =-7840;
14569: waveform_sig_loopback =-8062;
14570: waveform_sig_loopback =-8187;
14571: waveform_sig_loopback =-5499;
14572: waveform_sig_loopback =-6522;
14573: waveform_sig_loopback =-8902;
14574: waveform_sig_loopback =-6643;
14575: waveform_sig_loopback =-7264;
14576: waveform_sig_loopback =-7106;
14577: waveform_sig_loopback =-6805;
14578: waveform_sig_loopback =-8600;
14579: waveform_sig_loopback =-5715;
14580: waveform_sig_loopback =-7626;
14581: waveform_sig_loopback =-7682;
14582: waveform_sig_loopback =-6699;
14583: waveform_sig_loopback =-7310;
14584: waveform_sig_loopback =-7413;
14585: waveform_sig_loopback =-7217;
14586: waveform_sig_loopback =-6292;
14587: waveform_sig_loopback =-8413;
14588: waveform_sig_loopback =-6614;
14589: waveform_sig_loopback =-6903;
14590: waveform_sig_loopback =-7354;
14591: waveform_sig_loopback =-7669;
14592: waveform_sig_loopback =-6436;
14593: waveform_sig_loopback =-6714;
14594: waveform_sig_loopback =-8771;
14595: waveform_sig_loopback =-5844;
14596: waveform_sig_loopback =-6422;
14597: waveform_sig_loopback =-8858;
14598: waveform_sig_loopback =-6488;
14599: waveform_sig_loopback =-5998;
14600: waveform_sig_loopback =-7734;
14601: waveform_sig_loopback =-8026;
14602: waveform_sig_loopback =-5866;
14603: waveform_sig_loopback =-6899;
14604: waveform_sig_loopback =-7543;
14605: waveform_sig_loopback =-5513;
14606: waveform_sig_loopback =-10285;
14607: waveform_sig_loopback =-6031;
14608: waveform_sig_loopback =-4983;
14609: waveform_sig_loopback =-7778;
14610: waveform_sig_loopback =-7967;
14611: waveform_sig_loopback =-7482;
14612: waveform_sig_loopback =-5483;
14613: waveform_sig_loopback =-6242;
14614: waveform_sig_loopback =-8486;
14615: waveform_sig_loopback =-6382;
14616: waveform_sig_loopback =-6901;
14617: waveform_sig_loopback =-6711;
14618: waveform_sig_loopback =-6586;
14619: waveform_sig_loopback =-8054;
14620: waveform_sig_loopback =-5288;
14621: waveform_sig_loopback =-7490;
14622: waveform_sig_loopback =-7013;
14623: waveform_sig_loopback =-6248;
14624: waveform_sig_loopback =-7103;
14625: waveform_sig_loopback =-6652;
14626: waveform_sig_loopback =-6957;
14627: waveform_sig_loopback =-5818;
14628: waveform_sig_loopback =-7650;
14629: waveform_sig_loopback =-6633;
14630: waveform_sig_loopback =-5866;
14631: waveform_sig_loopback =-7131;
14632: waveform_sig_loopback =-7272;
14633: waveform_sig_loopback =-5334;
14634: waveform_sig_loopback =-6939;
14635: waveform_sig_loopback =-7755;
14636: waveform_sig_loopback =-5295;
14637: waveform_sig_loopback =-6267;
14638: waveform_sig_loopback =-7831;
14639: waveform_sig_loopback =-6207;
14640: waveform_sig_loopback =-5388;
14641: waveform_sig_loopback =-6992;
14642: waveform_sig_loopback =-7577;
14643: waveform_sig_loopback =-4979;
14644: waveform_sig_loopback =-6413;
14645: waveform_sig_loopback =-6845;
14646: waveform_sig_loopback =-4759;
14647: waveform_sig_loopback =-9744;
14648: waveform_sig_loopback =-5196;
14649: waveform_sig_loopback =-4146;
14650: waveform_sig_loopback =-7264;
14651: waveform_sig_loopback =-7242;
14652: waveform_sig_loopback =-6459;
14653: waveform_sig_loopback =-4873;
14654: waveform_sig_loopback =-5450;
14655: waveform_sig_loopback =-7637;
14656: waveform_sig_loopback =-5708;
14657: waveform_sig_loopback =-5862;
14658: waveform_sig_loopback =-5918;
14659: waveform_sig_loopback =-6004;
14660: waveform_sig_loopback =-6786;
14661: waveform_sig_loopback =-4706;
14662: waveform_sig_loopback =-6604;
14663: waveform_sig_loopback =-5868;
14664: waveform_sig_loopback =-5798;
14665: waveform_sig_loopback =-5788;
14666: waveform_sig_loopback =-5965;
14667: waveform_sig_loopback =-6169;
14668: waveform_sig_loopback =-4502;
14669: waveform_sig_loopback =-7152;
14670: waveform_sig_loopback =-5398;
14671: waveform_sig_loopback =-4830;
14672: waveform_sig_loopback =-6576;
14673: waveform_sig_loopback =-5803;
14674: waveform_sig_loopback =-4532;
14675: waveform_sig_loopback =-6163;
14676: waveform_sig_loopback =-6252;
14677: waveform_sig_loopback =-4515;
14678: waveform_sig_loopback =-5204;
14679: waveform_sig_loopback =-6717;
14680: waveform_sig_loopback =-5191;
14681: waveform_sig_loopback =-4098;
14682: waveform_sig_loopback =-6060;
14683: waveform_sig_loopback =-6539;
14684: waveform_sig_loopback =-3568;
14685: waveform_sig_loopback =-5575;
14686: waveform_sig_loopback =-5548;
14687: waveform_sig_loopback =-3608;
14688: waveform_sig_loopback =-8817;
14689: waveform_sig_loopback =-3689;
14690: waveform_sig_loopback =-2999;
14691: waveform_sig_loopback =-6371;
14692: waveform_sig_loopback =-5785;
14693: waveform_sig_loopback =-5329;
14694: waveform_sig_loopback =-3809;
14695: waveform_sig_loopback =-3970;
14696: waveform_sig_loopback =-6739;
14697: waveform_sig_loopback =-4293;
14698: waveform_sig_loopback =-4503;
14699: waveform_sig_loopback =-4968;
14700: waveform_sig_loopback =-4479;
14701: waveform_sig_loopback =-5596;
14702: waveform_sig_loopback =-3572;
14703: waveform_sig_loopback =-5006;
14704: waveform_sig_loopback =-4884;
14705: waveform_sig_loopback =-4433;
14706: waveform_sig_loopback =-4236;
14707: waveform_sig_loopback =-5084;
14708: waveform_sig_loopback =-4406;
14709: waveform_sig_loopback =-3376;
14710: waveform_sig_loopback =-5960;
14711: waveform_sig_loopback =-3606;
14712: waveform_sig_loopback =-3835;
14713: waveform_sig_loopback =-5080;
14714: waveform_sig_loopback =-4259;
14715: waveform_sig_loopback =-3362;
14716: waveform_sig_loopback =-4594;
14717: waveform_sig_loopback =-4889;
14718: waveform_sig_loopback =-3165;
14719: waveform_sig_loopback =-3662;
14720: waveform_sig_loopback =-5303;
14721: waveform_sig_loopback =-3863;
14722: waveform_sig_loopback =-2432;
14723: waveform_sig_loopback =-4904;
14724: waveform_sig_loopback =-5012;
14725: waveform_sig_loopback =-1762;
14726: waveform_sig_loopback =-4646;
14727: waveform_sig_loopback =-3587;
14728: waveform_sig_loopback =-2304;
14729: waveform_sig_loopback =-7616;
14730: waveform_sig_loopback =-1427;
14731: waveform_sig_loopback =-2232;
14732: waveform_sig_loopback =-4698;
14733: waveform_sig_loopback =-4045;
14734: waveform_sig_loopback =-4153;
14735: waveform_sig_loopback =-1821;
14736: waveform_sig_loopback =-2972;
14737: waveform_sig_loopback =-5090;
14738: waveform_sig_loopback =-2343;
14739: waveform_sig_loopback =-3412;
14740: waveform_sig_loopback =-3419;
14741: waveform_sig_loopback =-2748;
14742: waveform_sig_loopback =-4073;
14743: waveform_sig_loopback =-1883;
14744: waveform_sig_loopback =-3600;
14745: waveform_sig_loopback =-3369;
14746: waveform_sig_loopback =-2442;
14747: waveform_sig_loopback =-2875;
14748: waveform_sig_loopback =-3654;
14749: waveform_sig_loopback =-2360;
14750: waveform_sig_loopback =-2066;
14751: waveform_sig_loopback =-4294;
14752: waveform_sig_loopback =-1824;
14753: waveform_sig_loopback =-2546;
14754: waveform_sig_loopback =-3086;
14755: waveform_sig_loopback =-2742;
14756: waveform_sig_loopback =-1918;
14757: waveform_sig_loopback =-2546;
14758: waveform_sig_loopback =-3529;
14759: waveform_sig_loopback =-1341;
14760: waveform_sig_loopback =-1973;
14761: waveform_sig_loopback =-3912;
14762: waveform_sig_loopback =-1706;
14763: waveform_sig_loopback =-960;
14764: waveform_sig_loopback =-3421;
14765: waveform_sig_loopback =-2875;
14766: waveform_sig_loopback =-254;
14767: waveform_sig_loopback =-3079;
14768: waveform_sig_loopback =-1468;
14769: waveform_sig_loopback =-1094;
14770: waveform_sig_loopback =-5615;
14771: waveform_sig_loopback =492;
14772: waveform_sig_loopback =-915;
14773: waveform_sig_loopback =-2516;
14774: waveform_sig_loopback =-2602;
14775: waveform_sig_loopback =-2389;
14776: waveform_sig_loopback =360;
14777: waveform_sig_loopback =-1518;
14778: waveform_sig_loopback =-3246;
14779: waveform_sig_loopback =-534;
14780: waveform_sig_loopback =-1869;
14781: waveform_sig_loopback =-1023;
14782: waveform_sig_loopback =-1388;
14783: waveform_sig_loopback =-2448;
14784: waveform_sig_loopback =332;
14785: waveform_sig_loopback =-2080;
14786: waveform_sig_loopback =-1434;
14787: waveform_sig_loopback =-718;
14788: waveform_sig_loopback =-1234;
14789: waveform_sig_loopback =-1532;
14790: waveform_sig_loopback =-576;
14791: waveform_sig_loopback =-629;
14792: waveform_sig_loopback =-2011;
14793: waveform_sig_loopback =-127;
14794: waveform_sig_loopback =-811;
14795: waveform_sig_loopback =-1057;
14796: waveform_sig_loopback =-1184;
14797: waveform_sig_loopback =353;
14798: waveform_sig_loopback =-994;
14799: waveform_sig_loopback =-1835;
14800: waveform_sig_loopback =990;
14801: waveform_sig_loopback =-480;
14802: waveform_sig_loopback =-2022;
14803: waveform_sig_loopback =364;
14804: waveform_sig_loopback =673;
14805: waveform_sig_loopback =-1442;
14806: waveform_sig_loopback =-922;
14807: waveform_sig_loopback =1393;
14808: waveform_sig_loopback =-1039;
14809: waveform_sig_loopback =517;
14810: waveform_sig_loopback =339;
14811: waveform_sig_loopback =-3372;
14812: waveform_sig_loopback =2287;
14813: waveform_sig_loopback =922;
14814: waveform_sig_loopback =-516;
14815: waveform_sig_loopback =-1107;
14816: waveform_sig_loopback =-33;
14817: waveform_sig_loopback =2091;
14818: waveform_sig_loopback =39;
14819: waveform_sig_loopback =-966;
14820: waveform_sig_loopback =1122;
14821: waveform_sig_loopback =40;
14822: waveform_sig_loopback =1058;
14823: waveform_sig_loopback =126;
14824: waveform_sig_loopback =-169;
14825: waveform_sig_loopback =2124;
14826: waveform_sig_loopback =-460;
14827: waveform_sig_loopback =848;
14828: waveform_sig_loopback =965;
14829: waveform_sig_loopback =643;
14830: waveform_sig_loopback =562;
14831: waveform_sig_loopback =1090;
14832: waveform_sig_loopback =1421;
14833: waveform_sig_loopback =-53;
14834: waveform_sig_loopback =1496;
14835: waveform_sig_loopback =1425;
14836: waveform_sig_loopback =609;
14837: waveform_sig_loopback =743;
14838: waveform_sig_loopback =2482;
14839: waveform_sig_loopback =502;
14840: waveform_sig_loopback =405;
14841: waveform_sig_loopback =2868;
14842: waveform_sig_loopback =1054;
14843: waveform_sig_loopback =123;
14844: waveform_sig_loopback =2297;
14845: waveform_sig_loopback =2335;
14846: waveform_sig_loopback =561;
14847: waveform_sig_loopback =892;
14848: waveform_sig_loopback =3303;
14849: waveform_sig_loopback =943;
14850: waveform_sig_loopback =2154;
14851: waveform_sig_loopback =2311;
14852: waveform_sig_loopback =-1382;
14853: waveform_sig_loopback =4006;
14854: waveform_sig_loopback =3079;
14855: waveform_sig_loopback =1019;
14856: waveform_sig_loopback =846;
14857: waveform_sig_loopback =2153;
14858: waveform_sig_loopback =3538;
14859: waveform_sig_loopback =2175;
14860: waveform_sig_loopback =845;
14861: waveform_sig_loopback =2792;
14862: waveform_sig_loopback =2208;
14863: waveform_sig_loopback =2625;
14864: waveform_sig_loopback =1971;
14865: waveform_sig_loopback =1916;
14866: waveform_sig_loopback =3627;
14867: waveform_sig_loopback =1562;
14868: waveform_sig_loopback =2741;
14869: waveform_sig_loopback =2560;
14870: waveform_sig_loopback =2707;
14871: waveform_sig_loopback =2247;
14872: waveform_sig_loopback =2951;
14873: waveform_sig_loopback =3340;
14874: waveform_sig_loopback =1551;
14875: waveform_sig_loopback =3424;
14876: waveform_sig_loopback =3394;
14877: waveform_sig_loopback =2044;
14878: waveform_sig_loopback =2824;
14879: waveform_sig_loopback =4266;
14880: waveform_sig_loopback =1907;
14881: waveform_sig_loopback =2693;
14882: waveform_sig_loopback =4367;
14883: waveform_sig_loopback =2781;
14884: waveform_sig_loopback =2220;
14885: waveform_sig_loopback =3695;
14886: waveform_sig_loopback =4393;
14887: waveform_sig_loopback =2170;
14888: waveform_sig_loopback =2553;
14889: waveform_sig_loopback =5393;
14890: waveform_sig_loopback =2229;
14891: waveform_sig_loopback =4152;
14892: waveform_sig_loopback =3992;
14893: waveform_sig_loopback =99;
14894: waveform_sig_loopback =6133;
14895: waveform_sig_loopback =4599;
14896: waveform_sig_loopback =2504;
14897: waveform_sig_loopback =2868;
14898: waveform_sig_loopback =3760;
14899: waveform_sig_loopback =5262;
14900: waveform_sig_loopback =3955;
14901: waveform_sig_loopback =2335;
14902: waveform_sig_loopback =4738;
14903: waveform_sig_loopback =3921;
14904: waveform_sig_loopback =4216;
14905: waveform_sig_loopback =3781;
14906: waveform_sig_loopback =3642;
14907: waveform_sig_loopback =5129;
14908: waveform_sig_loopback =3389;
14909: waveform_sig_loopback =4300;
14910: waveform_sig_loopback =4149;
14911: waveform_sig_loopback =4687;
14912: waveform_sig_loopback =3465;
14913: waveform_sig_loopback =4884;
14914: waveform_sig_loopback =5000;
14915: waveform_sig_loopback =2837;
14916: waveform_sig_loopback =5536;
14917: waveform_sig_loopback =4627;
14918: waveform_sig_loopback =3707;
14919: waveform_sig_loopback =4782;
14920: waveform_sig_loopback =5382;
14921: waveform_sig_loopback =3839;
14922: waveform_sig_loopback =4203;
14923: waveform_sig_loopback =5760;
14924: waveform_sig_loopback =4635;
14925: waveform_sig_loopback =3540;
14926: waveform_sig_loopback =5481;
14927: waveform_sig_loopback =6037;
14928: waveform_sig_loopback =3428;
14929: waveform_sig_loopback =4422;
14930: waveform_sig_loopback =6969;
14931: waveform_sig_loopback =3479;
14932: waveform_sig_loopback =6105;
14933: waveform_sig_loopback =5186;
14934: waveform_sig_loopback =1670;
14935: waveform_sig_loopback =8015;
14936: waveform_sig_loopback =5722;
14937: waveform_sig_loopback =4072;
14938: waveform_sig_loopback =4518;
14939: waveform_sig_loopback =5012;
14940: waveform_sig_loopback =6950;
14941: waveform_sig_loopback =5305;
14942: waveform_sig_loopback =3606;
14943: waveform_sig_loopback =6502;
14944: waveform_sig_loopback =5019;
14945: waveform_sig_loopback =5618;
14946: waveform_sig_loopback =5348;
14947: waveform_sig_loopback =4774;
14948: waveform_sig_loopback =6750;
14949: waveform_sig_loopback =4832;
14950: waveform_sig_loopback =5422;
14951: waveform_sig_loopback =5883;
14952: waveform_sig_loopback =5770;
14953: waveform_sig_loopback =4732;
14954: waveform_sig_loopback =6701;
14955: waveform_sig_loopback =5723;
14956: waveform_sig_loopback =4498;
14957: waveform_sig_loopback =7007;
14958: waveform_sig_loopback =5475;
14959: waveform_sig_loopback =5455;
14960: waveform_sig_loopback =5821;
14961: waveform_sig_loopback =6680;
14962: waveform_sig_loopback =5264;
14963: waveform_sig_loopback =5252;
14964: waveform_sig_loopback =7305;
14965: waveform_sig_loopback =5746;
14966: waveform_sig_loopback =4647;
14967: waveform_sig_loopback =6880;
14968: waveform_sig_loopback =7091;
14969: waveform_sig_loopback =4566;
14970: waveform_sig_loopback =5854;
14971: waveform_sig_loopback =8000;
14972: waveform_sig_loopback =4507;
14973: waveform_sig_loopback =7710;
14974: waveform_sig_loopback =5809;
14975: waveform_sig_loopback =3012;
14976: waveform_sig_loopback =9463;
14977: waveform_sig_loopback =6369;
14978: waveform_sig_loopback =5531;
14979: waveform_sig_loopback =5483;
14980: waveform_sig_loopback =5998;
14981: waveform_sig_loopback =8465;
14982: waveform_sig_loopback =5852;
14983: waveform_sig_loopback =4929;
14984: waveform_sig_loopback =7814;
14985: waveform_sig_loopback =5556;
14986: waveform_sig_loopback =7246;
14987: waveform_sig_loopback =5990;
14988: waveform_sig_loopback =5821;
14989: waveform_sig_loopback =8131;
14990: waveform_sig_loopback =5211;
14991: waveform_sig_loopback =6815;
14992: waveform_sig_loopback =6820;
14993: waveform_sig_loopback =6455;
14994: waveform_sig_loopback =6135;
14995: waveform_sig_loopback =7291;
14996: waveform_sig_loopback =6706;
14997: waveform_sig_loopback =5648;
14998: waveform_sig_loopback =7642;
14999: waveform_sig_loopback =6589;
15000: waveform_sig_loopback =6191;
15001: waveform_sig_loopback =6784;
15002: waveform_sig_loopback =7499;
15003: waveform_sig_loopback =6123;
15004: waveform_sig_loopback =6085;
15005: waveform_sig_loopback =8222;
15006: waveform_sig_loopback =6577;
15007: waveform_sig_loopback =5234;
15008: waveform_sig_loopback =8241;
15009: waveform_sig_loopback =7489;
15010: waveform_sig_loopback =5297;
15011: waveform_sig_loopback =7102;
15012: waveform_sig_loopback =8188;
15013: waveform_sig_loopback =5748;
15014: waveform_sig_loopback =8408;
15015: waveform_sig_loopback =6107;
15016: waveform_sig_loopback =4460;
15017: waveform_sig_loopback =9673;
15018: waveform_sig_loopback =7237;
15019: waveform_sig_loopback =6392;
15020: waveform_sig_loopback =5664;
15021: waveform_sig_loopback =7307;
15022: waveform_sig_loopback =8879;
15023: waveform_sig_loopback =6268;
15024: waveform_sig_loopback =6053;
15025: waveform_sig_loopback =7944;
15026: waveform_sig_loopback =6482;
15027: waveform_sig_loopback =7970;
15028: waveform_sig_loopback =6152;
15029: waveform_sig_loopback =6951;
15030: waveform_sig_loopback =8459;
15031: waveform_sig_loopback =5816;
15032: waveform_sig_loopback =7614;
15033: waveform_sig_loopback =7021;
15034: waveform_sig_loopback =7237;
15035: waveform_sig_loopback =6680;
15036: waveform_sig_loopback =7812;
15037: waveform_sig_loopback =7141;
15038: waveform_sig_loopback =6273;
15039: waveform_sig_loopback =8127;
15040: waveform_sig_loopback =7059;
15041: waveform_sig_loopback =6767;
15042: waveform_sig_loopback =7010;
15043: waveform_sig_loopback =8339;
15044: waveform_sig_loopback =6258;
15045: waveform_sig_loopback =6519;
15046: waveform_sig_loopback =9037;
15047: waveform_sig_loopback =6319;
15048: waveform_sig_loopback =6110;
15049: waveform_sig_loopback =8600;
15050: waveform_sig_loopback =7454;
15051: waveform_sig_loopback =6229;
15052: waveform_sig_loopback =6997;
15053: waveform_sig_loopback =8685;
15054: waveform_sig_loopback =6221;
15055: waveform_sig_loopback =8311;
15056: waveform_sig_loopback =6635;
15057: waveform_sig_loopback =4670;
15058: waveform_sig_loopback =9947;
15059: waveform_sig_loopback =7765;
15060: waveform_sig_loopback =6120;
15061: waveform_sig_loopback =6238;
15062: waveform_sig_loopback =7665;
15063: waveform_sig_loopback =8729;
15064: waveform_sig_loopback =6774;
15065: waveform_sig_loopback =6120;
15066: waveform_sig_loopback =8086;
15067: waveform_sig_loopback =6792;
15068: waveform_sig_loopback =7943;
15069: waveform_sig_loopback =6369;
15070: waveform_sig_loopback =7228;
15071: waveform_sig_loopback =8299;
15072: waveform_sig_loopback =6041;
15073: waveform_sig_loopback =7816;
15074: waveform_sig_loopback =7048;
15075: waveform_sig_loopback =7322;
15076: waveform_sig_loopback =6749;
15077: waveform_sig_loopback =7752;
15078: waveform_sig_loopback =7309;
15079: waveform_sig_loopback =6214;
15080: waveform_sig_loopback =7911;
15081: waveform_sig_loopback =7504;
15082: waveform_sig_loopback =6174;
15083: waveform_sig_loopback =7426;
15084: waveform_sig_loopback =8055;
15085: waveform_sig_loopback =5757;
15086: waveform_sig_loopback =7295;
15087: waveform_sig_loopback =8314;
15088: waveform_sig_loopback =6183;
15089: waveform_sig_loopback =6274;
15090: waveform_sig_loopback =8209;
15091: waveform_sig_loopback =7662;
15092: waveform_sig_loopback =5662;
15093: waveform_sig_loopback =6782;
15094: waveform_sig_loopback =9030;
15095: waveform_sig_loopback =5485;
15096: waveform_sig_loopback =8418;
15097: waveform_sig_loopback =6260;
15098: waveform_sig_loopback =4351;
15099: waveform_sig_loopback =10155;
15100: waveform_sig_loopback =6990;
15101: waveform_sig_loopback =5916;
15102: waveform_sig_loopback =6268;
15103: waveform_sig_loopback =7203;
15104: waveform_sig_loopback =8417;
15105: waveform_sig_loopback =6359;
15106: waveform_sig_loopback =5914;
15107: waveform_sig_loopback =7722;
15108: waveform_sig_loopback =6451;
15109: waveform_sig_loopback =7405;
15110: waveform_sig_loopback =6160;
15111: waveform_sig_loopback =6931;
15112: waveform_sig_loopback =7519;
15113: waveform_sig_loopback =5965;
15114: waveform_sig_loopback =7162;
15115: waveform_sig_loopback =6531;
15116: waveform_sig_loopback =7125;
15117: waveform_sig_loopback =5807;
15118: waveform_sig_loopback =7675;
15119: waveform_sig_loopback =6718;
15120: waveform_sig_loopback =5401;
15121: waveform_sig_loopback =7949;
15122: waveform_sig_loopback =6458;
15123: waveform_sig_loopback =5818;
15124: waveform_sig_loopback =7135;
15125: waveform_sig_loopback =7121;
15126: waveform_sig_loopback =5662;
15127: waveform_sig_loopback =6426;
15128: waveform_sig_loopback =7648;
15129: waveform_sig_loopback =5987;
15130: waveform_sig_loopback =5447;
15131: waveform_sig_loopback =7572;
15132: waveform_sig_loopback =7030;
15133: waveform_sig_loopback =4944;
15134: waveform_sig_loopback =6513;
15135: waveform_sig_loopback =8048;
15136: waveform_sig_loopback =4637;
15137: waveform_sig_loopback =8235;
15138: waveform_sig_loopback =5077;
15139: waveform_sig_loopback =3762;
15140: waveform_sig_loopback =9663;
15141: waveform_sig_loopback =5988;
15142: waveform_sig_loopback =5238;
15143: waveform_sig_loopback =5468;
15144: waveform_sig_loopback =6363;
15145: waveform_sig_loopback =7889;
15146: waveform_sig_loopback =5376;
15147: waveform_sig_loopback =4977;
15148: waveform_sig_loopback =7205;
15149: waveform_sig_loopback =5492;
15150: waveform_sig_loopback =6563;
15151: waveform_sig_loopback =5383;
15152: waveform_sig_loopback =5881;
15153: waveform_sig_loopback =6915;
15154: waveform_sig_loopback =5093;
15155: waveform_sig_loopback =5980;
15156: waveform_sig_loopback =6071;
15157: waveform_sig_loopback =5995;
15158: waveform_sig_loopback =4913;
15159: waveform_sig_loopback =7069;
15160: waveform_sig_loopback =5256;
15161: waveform_sig_loopback =4932;
15162: waveform_sig_loopback =6904;
15163: waveform_sig_loopback =5203;
15164: waveform_sig_loopback =5250;
15165: waveform_sig_loopback =5890;
15166: waveform_sig_loopback =6217;
15167: waveform_sig_loopback =4733;
15168: waveform_sig_loopback =5266;
15169: waveform_sig_loopback =6816;
15170: waveform_sig_loopback =4816;
15171: waveform_sig_loopback =4324;
15172: waveform_sig_loopback =6748;
15173: waveform_sig_loopback =5783;
15174: waveform_sig_loopback =3758;
15175: waveform_sig_loopback =5752;
15176: waveform_sig_loopback =6657;
15177: waveform_sig_loopback =3631;
15178: waveform_sig_loopback =7345;
15179: waveform_sig_loopback =3456;
15180: waveform_sig_loopback =3127;
15181: waveform_sig_loopback =8486;
15182: waveform_sig_loopback =4586;
15183: waveform_sig_loopback =4384;
15184: waveform_sig_loopback =4083;
15185: waveform_sig_loopback =5278;
15186: waveform_sig_loopback =6931;
15187: waveform_sig_loopback =3733;
15188: waveform_sig_loopback =4092;
15189: waveform_sig_loopback =5997;
15190: waveform_sig_loopback =4025;
15191: waveform_sig_loopback =5734;
15192: waveform_sig_loopback =3783;
15193: waveform_sig_loopback =4776;
15194: waveform_sig_loopback =5837;
15195: waveform_sig_loopback =3422;
15196: waveform_sig_loopback =5017;
15197: waveform_sig_loopback =4745;
15198: waveform_sig_loopback =4407;
15199: waveform_sig_loopback =3912;
15200: waveform_sig_loopback =5574;
15201: waveform_sig_loopback =3846;
15202: waveform_sig_loopback =3903;
15203: waveform_sig_loopback =5222;
15204: waveform_sig_loopback =4037;
15205: waveform_sig_loopback =3934;
15206: waveform_sig_loopback =4355;
15207: waveform_sig_loopback =5028;
15208: waveform_sig_loopback =3158;
15209: waveform_sig_loopback =3927;
15210: waveform_sig_loopback =5542;
15211: waveform_sig_loopback =3149;
15212: waveform_sig_loopback =3041;
15213: waveform_sig_loopback =5535;
15214: waveform_sig_loopback =4011;
15215: waveform_sig_loopback =2483;
15216: waveform_sig_loopback =4481;
15217: waveform_sig_loopback =4871;
15218: waveform_sig_loopback =2500;
15219: waveform_sig_loopback =5713;
15220: waveform_sig_loopback =1700;
15221: waveform_sig_loopback =2165;
15222: waveform_sig_loopback =6587;
15223: waveform_sig_loopback =3224;
15224: waveform_sig_loopback =2910;
15225: waveform_sig_loopback =2286;
15226: waveform_sig_loopback =4191;
15227: waveform_sig_loopback =5137;
15228: waveform_sig_loopback =2051;
15229: waveform_sig_loopback =2896;
15230: waveform_sig_loopback =4088;
15231: waveform_sig_loopback =2649;
15232: waveform_sig_loopback =4242;
15233: waveform_sig_loopback =1860;
15234: waveform_sig_loopback =3593;
15235: waveform_sig_loopback =4006;
15236: waveform_sig_loopback =1760;
15237: waveform_sig_loopback =3695;
15238: waveform_sig_loopback =2850;
15239: waveform_sig_loopback =2893;
15240: waveform_sig_loopback =2472;
15241: waveform_sig_loopback =3668;
15242: waveform_sig_loopback =2337;
15243: waveform_sig_loopback =2341;
15244: waveform_sig_loopback =3356;
15245: waveform_sig_loopback =2700;
15246: waveform_sig_loopback =1987;
15247: waveform_sig_loopback =2816;
15248: waveform_sig_loopback =3529;
15249: waveform_sig_loopback =1056;
15250: waveform_sig_loopback =2689;
15251: waveform_sig_loopback =3696;
15252: waveform_sig_loopback =1244;
15253: waveform_sig_loopback =1700;
15254: waveform_sig_loopback =3582;
15255: waveform_sig_loopback =2328;
15256: waveform_sig_loopback =833;
15257: waveform_sig_loopback =2719;
15258: waveform_sig_loopback =3113;
15259: waveform_sig_loopback =861;
15260: waveform_sig_loopback =3929;
15261: waveform_sig_loopback =-163;
15262: waveform_sig_loopback =723;
15263: waveform_sig_loopback =4610;
15264: waveform_sig_loopback =1623;
15265: waveform_sig_loopback =938;
15266: waveform_sig_loopback =533;
15267: waveform_sig_loopback =2823;
15268: waveform_sig_loopback =2854;
15269: waveform_sig_loopback =541;
15270: waveform_sig_loopback =1162;
15271: waveform_sig_loopback =2011;
15272: waveform_sig_loopback =1282;
15273: waveform_sig_loopback =2071;
15274: waveform_sig_loopback =208;
15275: waveform_sig_loopback =2041;
15276: waveform_sig_loopback =1773;
15277: waveform_sig_loopback =307;
15278: waveform_sig_loopback =1798;
15279: waveform_sig_loopback =903;
15280: waveform_sig_loopback =1330;
15281: waveform_sig_loopback =450;
15282: waveform_sig_loopback =1971;
15283: waveform_sig_loopback =597;
15284: waveform_sig_loopback =302;
15285: waveform_sig_loopback =1753;
15286: waveform_sig_loopback =721;
15287: waveform_sig_loopback =95;
15288: waveform_sig_loopback =1175;
15289: waveform_sig_loopback =1475;
15290: waveform_sig_loopback =-816;
15291: waveform_sig_loopback =1057;
15292: waveform_sig_loopback =1686;
15293: waveform_sig_loopback =-738;
15294: waveform_sig_loopback =196;
15295: waveform_sig_loopback =1462;
15296: waveform_sig_loopback =594;
15297: waveform_sig_loopback =-1043;
15298: waveform_sig_loopback =772;
15299: waveform_sig_loopback =1504;
15300: waveform_sig_loopback =-1287;
15301: waveform_sig_loopback =2177;
15302: waveform_sig_loopback =-2132;
15303: waveform_sig_loopback =-1179;
15304: waveform_sig_loopback =2920;
15305: waveform_sig_loopback =-378;
15306: waveform_sig_loopback =-1154;
15307: waveform_sig_loopback =-1010;
15308: waveform_sig_loopback =794;
15309: waveform_sig_loopback =883;
15310: waveform_sig_loopback =-1182;
15311: waveform_sig_loopback =-980;
15312: waveform_sig_loopback =338;
15313: waveform_sig_loopback =-613;
15314: waveform_sig_loopback =-117;
15315: waveform_sig_loopback =-1366;
15316: waveform_sig_loopback =-5;
15317: waveform_sig_loopback =-205;
15318: waveform_sig_loopback =-1337;
15319: waveform_sig_loopback =-373;
15320: waveform_sig_loopback =-777;
15321: waveform_sig_loopback =-628;
15322: waveform_sig_loopback =-1575;
15323: waveform_sig_loopback =345;
15324: waveform_sig_loopback =-1568;
15325: waveform_sig_loopback =-1478;
15326: waveform_sig_loopback =-24;
15327: waveform_sig_loopback =-1294;
15328: waveform_sig_loopback =-1830;
15329: waveform_sig_loopback =-434;
15330: waveform_sig_loopback =-675;
15331: waveform_sig_loopback =-2596;
15332: waveform_sig_loopback =-619;
15333: waveform_sig_loopback =-571;
15334: waveform_sig_loopback =-2299;
15335: waveform_sig_loopback =-1884;
15336: waveform_sig_loopback =-421;
15337: waveform_sig_loopback =-1130;
15338: waveform_sig_loopback =-3290;
15339: waveform_sig_loopback =-742;
15340: waveform_sig_loopback =-503;
15341: waveform_sig_loopback =-3375;
15342: waveform_sig_loopback =642;
15343: waveform_sig_loopback =-4353;
15344: waveform_sig_loopback =-2858;
15345: waveform_sig_loopback =1265;
15346: waveform_sig_loopback =-2704;
15347: waveform_sig_loopback =-2791;
15348: waveform_sig_loopback =-2717;
15349: waveform_sig_loopback =-1406;
15350: waveform_sig_loopback =-600;
15351: waveform_sig_loopback =-3373;
15352: waveform_sig_loopback =-2722;
15353: waveform_sig_loopback =-1310;
15354: waveform_sig_loopback =-2810;
15355: waveform_sig_loopback =-1717;
15356: waveform_sig_loopback =-3290;
15357: waveform_sig_loopback =-1890;
15358: waveform_sig_loopback =-2013;
15359: waveform_sig_loopback =-3243;
15360: waveform_sig_loopback =-2222;
15361: waveform_sig_loopback =-2547;
15362: waveform_sig_loopback =-2553;
15363: waveform_sig_loopback =-3408;
15364: waveform_sig_loopback =-1335;
15365: waveform_sig_loopback =-3710;
15366: waveform_sig_loopback =-3208;
15367: waveform_sig_loopback =-1651;
15368: waveform_sig_loopback =-3558;
15369: waveform_sig_loopback =-3351;
15370: waveform_sig_loopback =-2260;
15371: waveform_sig_loopback =-2816;
15372: waveform_sig_loopback =-4022;
15373: waveform_sig_loopback =-2787;
15374: waveform_sig_loopback =-2186;
15375: waveform_sig_loopback =-4087;
15376: waveform_sig_loopback =-3999;
15377: waveform_sig_loopback =-1693;
15378: waveform_sig_loopback =-3336;
15379: waveform_sig_loopback =-4968;
15380: waveform_sig_loopback =-2217;
15381: waveform_sig_loopback =-2761;
15382: waveform_sig_loopback =-4767;
15383: waveform_sig_loopback =-1117;
15384: waveform_sig_loopback =-6436;
15385: waveform_sig_loopback =-4158;
15386: waveform_sig_loopback =-693;
15387: waveform_sig_loopback =-4471;
15388: waveform_sig_loopback =-4429;
15389: waveform_sig_loopback =-4621;
15390: waveform_sig_loopback =-2987;
15391: waveform_sig_loopback =-2230;
15392: waveform_sig_loopback =-5325;
15393: waveform_sig_loopback =-4268;
15394: waveform_sig_loopback =-3006;
15395: waveform_sig_loopback =-4652;
15396: waveform_sig_loopback =-3168;
15397: waveform_sig_loopback =-5143;
15398: waveform_sig_loopback =-3554;
15399: waveform_sig_loopback =-3500;
15400: waveform_sig_loopback =-5153;
15401: waveform_sig_loopback =-3796;
15402: waveform_sig_loopback =-4122;
15403: waveform_sig_loopback =-4518;
15404: waveform_sig_loopback =-4741;
15405: waveform_sig_loopback =-3078;
15406: waveform_sig_loopback =-5568;
15407: waveform_sig_loopback =-4353;
15408: waveform_sig_loopback =-3621;
15409: waveform_sig_loopback =-5053;
15410: waveform_sig_loopback =-4793;
15411: waveform_sig_loopback =-4111;
15412: waveform_sig_loopback =-4103;
15413: waveform_sig_loopback =-5792;
15414: waveform_sig_loopback =-4348;
15415: waveform_sig_loopback =-3493;
15416: waveform_sig_loopback =-6012;
15417: waveform_sig_loopback =-5331;
15418: waveform_sig_loopback =-3170;
15419: waveform_sig_loopback =-5152;
15420: waveform_sig_loopback =-6352;
15421: waveform_sig_loopback =-3636;
15422: waveform_sig_loopback =-4495;
15423: waveform_sig_loopback =-6049;
15424: waveform_sig_loopback =-2801;
15425: waveform_sig_loopback =-8183;
15426: waveform_sig_loopback =-5153;
15427: waveform_sig_loopback =-2423;
15428: waveform_sig_loopback =-6022;
15429: waveform_sig_loopback =-5710;
15430: waveform_sig_loopback =-6333;
15431: waveform_sig_loopback =-4135;
15432: waveform_sig_loopback =-3808;
15433: waveform_sig_loopback =-7131;
15434: waveform_sig_loopback =-5203;
15435: waveform_sig_loopback =-4964;
15436: waveform_sig_loopback =-5778;
15437: waveform_sig_loopback =-4426;
15438: waveform_sig_loopback =-7108;
15439: waveform_sig_loopback =-4586;
15440: waveform_sig_loopback =-4981;
15441: waveform_sig_loopback =-6561;
15442: waveform_sig_loopback =-4851;
15443: waveform_sig_loopback =-5930;
15444: waveform_sig_loopback =-5661;
15445: waveform_sig_loopback =-5789;
15446: waveform_sig_loopback =-4909;
15447: waveform_sig_loopback =-6623;
15448: waveform_sig_loopback =-5757;
15449: waveform_sig_loopback =-5054;
15450: waveform_sig_loopback =-6205;
15451: waveform_sig_loopback =-6425;
15452: waveform_sig_loopback =-5175;
15453: waveform_sig_loopback =-5447;
15454: waveform_sig_loopback =-7324;
15455: waveform_sig_loopback =-5449;
15456: waveform_sig_loopback =-4733;
15457: waveform_sig_loopback =-7449;
15458: waveform_sig_loopback =-6401;
15459: waveform_sig_loopback =-4415;
15460: waveform_sig_loopback =-6604;
15461: waveform_sig_loopback =-7305;
15462: waveform_sig_loopback =-5024;
15463: waveform_sig_loopback =-5858;
15464: waveform_sig_loopback =-6827;
15465: waveform_sig_loopback =-4401;
15466: waveform_sig_loopback =-9303;
15467: waveform_sig_loopback =-5977;
15468: waveform_sig_loopback =-4061;
15469: waveform_sig_loopback =-6753;
15470: waveform_sig_loopback =-7207;
15471: waveform_sig_loopback =-7430;
15472: waveform_sig_loopback =-4758;
15473: waveform_sig_loopback =-5547;
15474: waveform_sig_loopback =-7888;
15475: waveform_sig_loopback =-6224;
15476: waveform_sig_loopback =-6250;
15477: waveform_sig_loopback =-6431;
15478: waveform_sig_loopback =-6041;
15479: waveform_sig_loopback =-7869;
15480: waveform_sig_loopback =-5185;
15481: waveform_sig_loopback =-6738;
15482: waveform_sig_loopback =-7200;
15483: waveform_sig_loopback =-6025;
15484: waveform_sig_loopback =-6821;
15485: waveform_sig_loopback =-6592;
15486: waveform_sig_loopback =-7055;
15487: waveform_sig_loopback =-5591;
15488: waveform_sig_loopback =-7699;
15489: waveform_sig_loopback =-6617;
15490: waveform_sig_loopback =-6106;
15491: waveform_sig_loopback =-6980;
15492: waveform_sig_loopback =-7357;
15493: waveform_sig_loopback =-6089;
15494: waveform_sig_loopback =-6194;
15495: waveform_sig_loopback =-8427;
15496: waveform_sig_loopback =-5845;
15497: waveform_sig_loopback =-5913;
15498: waveform_sig_loopback =-8503;
15499: waveform_sig_loopback =-6569;
15500: waveform_sig_loopback =-5762;
15501: waveform_sig_loopback =-7211;
15502: waveform_sig_loopback =-8009;
15503: waveform_sig_loopback =-6056;
15504: waveform_sig_loopback =-6182;
15505: waveform_sig_loopback =-7999;
15506: waveform_sig_loopback =-5096;
15507: waveform_sig_loopback =-9843;
15508: waveform_sig_loopback =-6996;
15509: waveform_sig_loopback =-4388;
15510: waveform_sig_loopback =-7725;
15511: waveform_sig_loopback =-8089;
15512: waveform_sig_loopback =-7542;
15513: waveform_sig_loopback =-5919;
15514: waveform_sig_loopback =-6035;
15515: waveform_sig_loopback =-8389;
15516: waveform_sig_loopback =-7087;
15517: waveform_sig_loopback =-6628;
15518: waveform_sig_loopback =-7154;
15519: waveform_sig_loopback =-6719;
15520: waveform_sig_loopback =-8159;
15521: waveform_sig_loopback =-5992;
15522: waveform_sig_loopback =-7298;
15523: waveform_sig_loopback =-7594;
15524: waveform_sig_loopback =-6696;
15525: waveform_sig_loopback =-7325;
15526: waveform_sig_loopback =-7114;
15527: waveform_sig_loopback =-7577;
15528: waveform_sig_loopback =-6123;
15529: waveform_sig_loopback =-8064;
15530: waveform_sig_loopback =-7365;
15531: waveform_sig_loopback =-6266;
15532: waveform_sig_loopback =-7583;
15533: waveform_sig_loopback =-7970;
15534: waveform_sig_loopback =-5985;
15535: waveform_sig_loopback =-7316;
15536: waveform_sig_loopback =-8449;
15537: waveform_sig_loopback =-6090;
15538: waveform_sig_loopback =-6825;
15539: waveform_sig_loopback =-8321;
15540: waveform_sig_loopback =-7262;
15541: waveform_sig_loopback =-6087;
15542: waveform_sig_loopback =-7355;
15543: waveform_sig_loopback =-8776;
15544: waveform_sig_loopback =-5851;
15545: waveform_sig_loopback =-6763;
15546: waveform_sig_loopback =-8408;
15547: waveform_sig_loopback =-4995;
15548: waveform_sig_loopback =-10624;
15549: waveform_sig_loopback =-6867;
15550: waveform_sig_loopback =-4556;
15551: waveform_sig_loopback =-8426;
15552: waveform_sig_loopback =-7968;
15553: waveform_sig_loopback =-7778;
15554: waveform_sig_loopback =-6241;
15555: waveform_sig_loopback =-6067;
15556: waveform_sig_loopback =-8815;
15557: waveform_sig_loopback =-7049;
15558: waveform_sig_loopback =-6770;
15559: waveform_sig_loopback =-7427;
15560: waveform_sig_loopback =-6850;
15561: waveform_sig_loopback =-8177;
15562: waveform_sig_loopback =-6188;
15563: waveform_sig_loopback =-7500;
15564: waveform_sig_loopback =-7473;
15565: waveform_sig_loopback =-7034;
15566: waveform_sig_loopback =-7156;
15567: waveform_sig_loopback =-7197;
15568: waveform_sig_loopback =-7839;
15569: waveform_sig_loopback =-5681;
15570: waveform_sig_loopback =-8560;
15571: waveform_sig_loopback =-7116;
15572: waveform_sig_loopback =-6014;
15573: waveform_sig_loopback =-8177;
15574: waveform_sig_loopback =-7244;
15575: waveform_sig_loopback =-6266;
15576: waveform_sig_loopback =-7446;
15577: waveform_sig_loopback =-7803;
15578: waveform_sig_loopback =-6599;
15579: waveform_sig_loopback =-6321;
15580: waveform_sig_loopback =-8395;
15581: waveform_sig_loopback =-7241;
15582: waveform_sig_loopback =-5492;
15583: waveform_sig_loopback =-7767;
15584: waveform_sig_loopback =-8360;
15585: waveform_sig_loopback =-5495;
15586: waveform_sig_loopback =-6996;
15587: waveform_sig_loopback =-7830;
15588: waveform_sig_loopback =-4996;
15589: waveform_sig_loopback =-10519;
15590: waveform_sig_loopback =-6271;
15591: waveform_sig_loopback =-4562;
15592: waveform_sig_loopback =-8180;
15593: waveform_sig_loopback =-7632;
15594: waveform_sig_loopback =-7612;
15595: waveform_sig_loopback =-5858;
15596: waveform_sig_loopback =-5664;
15597: waveform_sig_loopback =-8779;
15598: waveform_sig_loopback =-6583;
15599: waveform_sig_loopback =-6405;
15600: waveform_sig_loopback =-7257;
15601: waveform_sig_loopback =-6261;
15602: waveform_sig_loopback =-7947;
15603: waveform_sig_loopback =-5828;
15604: waveform_sig_loopback =-6819;
15605: waveform_sig_loopback =-7360;
15606: waveform_sig_loopback =-6531;
15607: waveform_sig_loopback =-6465;
15608: waveform_sig_loopback =-7243;
15609: waveform_sig_loopback =-6794;
15610: waveform_sig_loopback =-5499;
15611: waveform_sig_loopback =-8292;
15612: waveform_sig_loopback =-5962;
15613: waveform_sig_loopback =-6210;
15614: waveform_sig_loopback =-7257;
15615: waveform_sig_loopback =-6726;
15616: waveform_sig_loopback =-6010;
15617: waveform_sig_loopback =-6466;
15618: waveform_sig_loopback =-7684;
15619: waveform_sig_loopback =-5766;
15620: waveform_sig_loopback =-5717;
15621: waveform_sig_loopback =-8004;
15622: waveform_sig_loopback =-6463;
15623: waveform_sig_loopback =-4876;
15624: waveform_sig_loopback =-7244;
15625: waveform_sig_loopback =-7652;
15626: waveform_sig_loopback =-4702;
15627: waveform_sig_loopback =-6673;
15628: waveform_sig_loopback =-6726;
15629: waveform_sig_loopback =-4545;
15630: waveform_sig_loopback =-10092;
15631: waveform_sig_loopback =-4899;
15632: waveform_sig_loopback =-4300;
15633: waveform_sig_loopback =-7320;
15634: waveform_sig_loopback =-6787;
15635: waveform_sig_loopback =-7071;
15636: waveform_sig_loopback =-4675;
15637: waveform_sig_loopback =-5189;
15638: waveform_sig_loopback =-8141;
15639: waveform_sig_loopback =-5354;
15640: waveform_sig_loopback =-5968;
15641: waveform_sig_loopback =-6300;
15642: waveform_sig_loopback =-5389;
15643: waveform_sig_loopback =-7411;
15644: waveform_sig_loopback =-4677;
15645: waveform_sig_loopback =-6135;
15646: waveform_sig_loopback =-6679;
15647: waveform_sig_loopback =-5254;
15648: waveform_sig_loopback =-5947;
15649: waveform_sig_loopback =-6335;
15650: waveform_sig_loopback =-5556;
15651: waveform_sig_loopback =-5093;
15652: waveform_sig_loopback =-6952;
15653: waveform_sig_loopback =-5150;
15654: waveform_sig_loopback =-5438;
15655: waveform_sig_loopback =-5920;
15656: waveform_sig_loopback =-6122;
15657: waveform_sig_loopback =-4791;
15658: waveform_sig_loopback =-5497;
15659: waveform_sig_loopback =-6864;
15660: waveform_sig_loopback =-4409;
15661: waveform_sig_loopback =-4966;
15662: waveform_sig_loopback =-7000;
15663: waveform_sig_loopback =-5180;
15664: waveform_sig_loopback =-3951;
15665: waveform_sig_loopback =-6293;
15666: waveform_sig_loopback =-6413;
15667: waveform_sig_loopback =-3623;
15668: waveform_sig_loopback =-5764;
15669: waveform_sig_loopback =-5250;
15670: waveform_sig_loopback =-3854;
15671: waveform_sig_loopback =-8825;
15672: waveform_sig_loopback =-3482;
15673: waveform_sig_loopback =-3629;
15674: waveform_sig_loopback =-5747;
15675: waveform_sig_loopback =-5931;
15676: waveform_sig_loopback =-5831;
15677: waveform_sig_loopback =-3118;
15678: waveform_sig_loopback =-4590;
15679: waveform_sig_loopback =-6504;
15680: waveform_sig_loopback =-4120;
15681: waveform_sig_loopback =-5048;
15682: waveform_sig_loopback =-4508;
15683: waveform_sig_loopback =-4561;
15684: waveform_sig_loopback =-5914;
15685: waveform_sig_loopback =-3086;
15686: waveform_sig_loopback =-5355;
15687: waveform_sig_loopback =-4904;
15688: waveform_sig_loopback =-4079;
15689: waveform_sig_loopback =-4763;
15690: waveform_sig_loopback =-4675;
15691: waveform_sig_loopback =-4446;
15692: waveform_sig_loopback =-3688;
15693: waveform_sig_loopback =-5493;
15694: waveform_sig_loopback =-3974;
15695: waveform_sig_loopback =-3891;
15696: waveform_sig_loopback =-4614;
15697: waveform_sig_loopback =-4927;
15698: waveform_sig_loopback =-3136;
15699: waveform_sig_loopback =-4340;
15700: waveform_sig_loopback =-5484;
15701: waveform_sig_loopback =-2740;
15702: waveform_sig_loopback =-3896;
15703: waveform_sig_loopback =-5451;
15704: waveform_sig_loopback =-3591;
15705: waveform_sig_loopback =-2870;
15706: waveform_sig_loopback =-4696;
15707: waveform_sig_loopback =-4908;
15708: waveform_sig_loopback =-2275;
15709: waveform_sig_loopback =-4206;
15710: waveform_sig_loopback =-3787;
15711: waveform_sig_loopback =-2553;
15712: waveform_sig_loopback =-7096;
15713: waveform_sig_loopback =-2053;
15714: waveform_sig_loopback =-2081;
15715: waveform_sig_loopback =-4193;
15716: waveform_sig_loopback =-4697;
15717: waveform_sig_loopback =-3774;
15718: waveform_sig_loopback =-1839;
15719: waveform_sig_loopback =-3136;
15720: waveform_sig_loopback =-4644;
15721: waveform_sig_loopback =-2923;
15722: waveform_sig_loopback =-3224;
15723: waveform_sig_loopback =-2926;
15724: waveform_sig_loopback =-3339;
15725: waveform_sig_loopback =-3945;
15726: waveform_sig_loopback =-1747;
15727: waveform_sig_loopback =-3781;
15728: waveform_sig_loopback =-3031;
15729: waveform_sig_loopback =-2864;
15730: waveform_sig_loopback =-2865;
15731: waveform_sig_loopback =-3098;
15732: waveform_sig_loopback =-2958;
15733: waveform_sig_loopback =-1835;
15734: waveform_sig_loopback =-4026;
15735: waveform_sig_loopback =-2334;
15736: waveform_sig_loopback =-2042;
15737: waveform_sig_loopback =-3245;
15738: waveform_sig_loopback =-2990;
15739: waveform_sig_loopback =-1474;
15740: waveform_sig_loopback =-2912;
15741: waveform_sig_loopback =-3425;
15742: waveform_sig_loopback =-1170;
15743: waveform_sig_loopback =-2263;
15744: waveform_sig_loopback =-3589;
15745: waveform_sig_loopback =-1799;
15746: waveform_sig_loopback =-1207;
15747: waveform_sig_loopback =-2886;
15748: waveform_sig_loopback =-3210;
15749: waveform_sig_loopback =-462;
15750: waveform_sig_loopback =-2434;
15751: waveform_sig_loopback =-2192;
15752: waveform_sig_loopback =-600;
15753: waveform_sig_loopback =-5430;
15754: waveform_sig_loopback =-252;
15755: waveform_sig_loopback =-13;
15756: waveform_sig_loopback =-2918;
15757: waveform_sig_loopback =-2710;
15758: waveform_sig_loopback =-1805;
15759: waveform_sig_loopback =-455;
15760: waveform_sig_loopback =-953;
15761: waveform_sig_loopback =-3160;
15762: waveform_sig_loopback =-1048;
15763: waveform_sig_loopback =-1202;
15764: waveform_sig_loopback =-1526;
15765: waveform_sig_loopback =-1243;
15766: waveform_sig_loopback =-2152;
15767: waveform_sig_loopback =-194;
15768: waveform_sig_loopback =-1705;
15769: waveform_sig_loopback =-1445;
15770: waveform_sig_loopback =-968;
15771: waveform_sig_loopback =-928;
15772: waveform_sig_loopback =-1568;
15773: waveform_sig_loopback =-904;
15774: waveform_sig_loopback =-84;
15775: waveform_sig_loopback =-2270;
15776: waveform_sig_loopback =-317;
15777: waveform_sig_loopback =-274;
15778: waveform_sig_loopback =-1489;
15779: waveform_sig_loopback =-990;
15780: waveform_sig_loopback =330;
15781: waveform_sig_loopback =-1208;
15782: waveform_sig_loopback =-1306;
15783: waveform_sig_loopback =562;
15784: waveform_sig_loopback =-634;
15785: waveform_sig_loopback =-1478;
15786: waveform_sig_loopback =-82;
15787: waveform_sig_loopback =875;
15788: waveform_sig_loopback =-1358;
15789: waveform_sig_loopback =-1487;
15790: waveform_sig_loopback =2098;
15791: waveform_sig_loopback =-1162;
15792: waveform_sig_loopback =-53;
15793: waveform_sig_loopback =1113;
15794: waveform_sig_loopback =-3800;
15795: waveform_sig_loopback =2268;
15796: waveform_sig_loopback =1291;
15797: waveform_sig_loopback =-1140;
15798: waveform_sig_loopback =-415;
15799: waveform_sig_loopback =-299;
15800: waveform_sig_loopback =1618;
15801: waveform_sig_loopback =833;
15802: waveform_sig_loopback =-1503;
15803: waveform_sig_loopback =1255;
15804: waveform_sig_loopback =264;
15805: waveform_sig_loopback =434;
15806: waveform_sig_loopback =855;
15807: waveform_sig_loopback =-534;
15808: waveform_sig_loopback =1893;
15809: waveform_sig_loopback =86;
15810: waveform_sig_loopback =439;
15811: waveform_sig_loopback =1008;
15812: waveform_sig_loopback =822;
15813: waveform_sig_loopback =309;
15814: waveform_sig_loopback =1126;
15815: waveform_sig_loopback =1709;
15816: waveform_sig_loopback =-512;
15817: waveform_sig_loopback =1825;
15818: waveform_sig_loopback =1447;
15819: waveform_sig_loopback =273;
15820: waveform_sig_loopback =1229;
15821: waveform_sig_loopback =1927;
15822: waveform_sig_loopback =815;
15823: waveform_sig_loopback =623;
15824: waveform_sig_loopback =2148;
15825: waveform_sig_loopback =1800;
15826: waveform_sig_loopback =-27;
15827: waveform_sig_loopback =1824;
15828: waveform_sig_loopback =2987;
15829: waveform_sig_loopback =160;
15830: waveform_sig_loopback =996;
15831: waveform_sig_loopback =3512;
15832: waveform_sig_loopback =427;
15833: waveform_sig_loopback =2615;
15834: waveform_sig_loopback =2314;
15835: waveform_sig_loopback =-1781;
15836: waveform_sig_loopback =4409;
15837: waveform_sig_loopback =2759;
15838: waveform_sig_loopback =1179;
15839: waveform_sig_loopback =1028;
15840: waveform_sig_loopback =1619;
15841: waveform_sig_loopback =3953;
15842: waveform_sig_loopback =2173;
15843: waveform_sig_loopback =533;
15844: waveform_sig_loopback =3169;
15845: waveform_sig_loopback =2004;
15846: waveform_sig_loopback =2575;
15847: waveform_sig_loopback =2329;
15848: waveform_sig_loopback =1406;
15849: waveform_sig_loopback =3869;
15850: waveform_sig_loopback =1822;
15851: waveform_sig_loopback =2232;
15852: waveform_sig_loopback =2918;
15853: waveform_sig_loopback =2712;
15854: waveform_sig_loopback =1931;
15855: waveform_sig_loopback =3327;
15856: waveform_sig_loopback =3083;
15857: waveform_sig_loopback =1536;
15858: waveform_sig_loopback =3822;
15859: waveform_sig_loopback =2728;
15860: waveform_sig_loopback =2683;
15861: waveform_sig_loopback =2632;
15862: waveform_sig_loopback =3832;
15863: waveform_sig_loopback =2833;
15864: waveform_sig_loopback =1931;
15865: waveform_sig_loopback =4536;
15866: waveform_sig_loopback =3211;
15867: waveform_sig_loopback =1624;
15868: waveform_sig_loopback =4127;
15869: waveform_sig_loopback =4232;
15870: waveform_sig_loopback =2066;
15871: waveform_sig_loopback =2886;
15872: waveform_sig_loopback =5036;
15873: waveform_sig_loopback =2418;
15874: waveform_sig_loopback =4332;
15875: waveform_sig_loopback =3845;
15876: waveform_sig_loopback =204;
15877: waveform_sig_loopback =6111;
15878: waveform_sig_loopback =4483;
15879: waveform_sig_loopback =2869;
15880: waveform_sig_loopback =2731;
15881: waveform_sig_loopback =3466;
15882: waveform_sig_loopback =5645;
15883: waveform_sig_loopback =3756;
15884: waveform_sig_loopback =2294;
15885: waveform_sig_loopback =5019;
15886: waveform_sig_loopback =3373;
15887: waveform_sig_loopback =4588;
15888: waveform_sig_loopback =3821;
15889: waveform_sig_loopback =3128;
15890: waveform_sig_loopback =5778;
15891: waveform_sig_loopback =3039;
15892: waveform_sig_loopback =4216;
15893: waveform_sig_loopback =4599;
15894: waveform_sig_loopback =4035;
15895: waveform_sig_loopback =3939;
15896: waveform_sig_loopback =4742;
15897: waveform_sig_loopback =4671;
15898: waveform_sig_loopback =3428;
15899: waveform_sig_loopback =4982;
15900: waveform_sig_loopback =4714;
15901: waveform_sig_loopback =4080;
15902: waveform_sig_loopback =4097;
15903: waveform_sig_loopback =5776;
15904: waveform_sig_loopback =3920;
15905: waveform_sig_loopback =3728;
15906: waveform_sig_loopback =6183;
15907: waveform_sig_loopback =4452;
15908: waveform_sig_loopback =3370;
15909: waveform_sig_loopback =5705;
15910: waveform_sig_loopback =5643;
15911: waveform_sig_loopback =3702;
15912: waveform_sig_loopback =4447;
15913: waveform_sig_loopback =6545;
15914: waveform_sig_loopback =4001;
15915: waveform_sig_loopback =5816;
15916: waveform_sig_loopback =5215;
15917: waveform_sig_loopback =1888;
15918: waveform_sig_loopback =7573;
15919: waveform_sig_loopback =5930;
15920: waveform_sig_loopback =4372;
15921: waveform_sig_loopback =4047;
15922: waveform_sig_loopback =5213;
15923: waveform_sig_loopback =7029;
15924: waveform_sig_loopback =4974;
15925: waveform_sig_loopback =4127;
15926: waveform_sig_loopback =6164;
15927: waveform_sig_loopback =4909;
15928: waveform_sig_loopback =6175;
15929: waveform_sig_loopback =4811;
15930: waveform_sig_loopback =5059;
15931: waveform_sig_loopback =6890;
15932: waveform_sig_loopback =4303;
15933: waveform_sig_loopback =6039;
15934: waveform_sig_loopback =5495;
15935: waveform_sig_loopback =5706;
15936: waveform_sig_loopback =5271;
15937: waveform_sig_loopback =5932;
15938: waveform_sig_loopback =6252;
15939: waveform_sig_loopback =4487;
15940: waveform_sig_loopback =6514;
15941: waveform_sig_loopback =6060;
15942: waveform_sig_loopback =5089;
15943: waveform_sig_loopback =5772;
15944: waveform_sig_loopback =6930;
15945: waveform_sig_loopback =5085;
15946: waveform_sig_loopback =5196;
15947: waveform_sig_loopback =7445;
15948: waveform_sig_loopback =5561;
15949: waveform_sig_loopback =4696;
15950: waveform_sig_loopback =7069;
15951: waveform_sig_loopback =6630;
15952: waveform_sig_loopback =5110;
15953: waveform_sig_loopback =5544;
15954: waveform_sig_loopback =7723;
15955: waveform_sig_loopback =5308;
15956: waveform_sig_loopback =6805;
15957: waveform_sig_loopback =6482;
15958: waveform_sig_loopback =3024;
15959: waveform_sig_loopback =8707;
15960: waveform_sig_loopback =7295;
15961: waveform_sig_loopback =5058;
15962: waveform_sig_loopback =5392;
15963: waveform_sig_loopback =6478;
15964: waveform_sig_loopback =7762;
15965: waveform_sig_loopback =6349;
15966: waveform_sig_loopback =4981;
15967: waveform_sig_loopback =7230;
15968: waveform_sig_loopback =6209;
15969: waveform_sig_loopback =6869;
15970: waveform_sig_loopback =5983;
15971: waveform_sig_loopback =6213;
15972: waveform_sig_loopback =7623;
15973: waveform_sig_loopback =5548;
15974: waveform_sig_loopback =6862;
15975: waveform_sig_loopback =6471;
15976: waveform_sig_loopback =6831;
15977: waveform_sig_loopback =6001;
15978: waveform_sig_loopback =7068;
15979: waveform_sig_loopback =7153;
15980: waveform_sig_loopback =5352;
15981: waveform_sig_loopback =7543;
15982: waveform_sig_loopback =7010;
15983: waveform_sig_loopback =5812;
15984: waveform_sig_loopback =6895;
15985: waveform_sig_loopback =7753;
15986: waveform_sig_loopback =5707;
15987: waveform_sig_loopback =6494;
15988: waveform_sig_loopback =8026;
15989: waveform_sig_loopback =6358;
15990: waveform_sig_loopback =5810;
15991: waveform_sig_loopback =7593;
15992: waveform_sig_loopback =7747;
15993: waveform_sig_loopback =5687;
15994: waveform_sig_loopback =6285;
15995: waveform_sig_loopback =8910;
15996: waveform_sig_loopback =5514;
15997: waveform_sig_loopback =7966;
15998: waveform_sig_loopback =7051;
15999: waveform_sig_loopback =3575;
16000: waveform_sig_loopback =9970;
16001: waveform_sig_loopback =7542;
16002: waveform_sig_loopback =5746;
16003: waveform_sig_loopback =6403;
16004: waveform_sig_loopback =6909;
16005: waveform_sig_loopback =8627;
16006: waveform_sig_loopback =6919;
16007: waveform_sig_loopback =5531;
16008: waveform_sig_loopback =8116;
16009: waveform_sig_loopback =6714;
16010: waveform_sig_loopback =7389;
16011: waveform_sig_loopback =6748;
16012: waveform_sig_loopback =6758;
16013: waveform_sig_loopback =8139;
16014: waveform_sig_loopback =6306;
16015: waveform_sig_loopback =7232;
16016: waveform_sig_loopback =7123;
16017: waveform_sig_loopback =7460;
16018: waveform_sig_loopback =6252;
16019: waveform_sig_loopback =7923;
16020: waveform_sig_loopback =7422;
16021: waveform_sig_loopback =5759;
16022: waveform_sig_loopback =8373;
16023: waveform_sig_loopback =7095;
16024: waveform_sig_loopback =6403;
16025: waveform_sig_loopback =7572;
16026: waveform_sig_loopback =7780;
16027: waveform_sig_loopback =6427;
16028: waveform_sig_loopback =6867;
16029: waveform_sig_loopback =8306;
16030: waveform_sig_loopback =6990;
16031: waveform_sig_loopback =5895;
16032: waveform_sig_loopback =8191;
16033: waveform_sig_loopback =8141;
16034: waveform_sig_loopback =5648;
16035: waveform_sig_loopback =7052;
16036: waveform_sig_loopback =9102;
16037: waveform_sig_loopback =5586;
16038: waveform_sig_loopback =8737;
16039: waveform_sig_loopback =6794;
16040: waveform_sig_loopback =4065;
16041: waveform_sig_loopback =10489;
16042: waveform_sig_loopback =7374;
16043: waveform_sig_loopback =6276;
16044: waveform_sig_loopback =6472;
16045: waveform_sig_loopback =7046;
16046: waveform_sig_loopback =9133;
16047: waveform_sig_loopback =6750;
16048: waveform_sig_loopback =5780;
16049: waveform_sig_loopback =8451;
16050: waveform_sig_loopback =6624;
16051: waveform_sig_loopback =7714;
16052: waveform_sig_loopback =6788;
16053: waveform_sig_loopback =6743;
16054: waveform_sig_loopback =8457;
16055: waveform_sig_loopback =6278;
16056: waveform_sig_loopback =7240;
16057: waveform_sig_loopback =7421;
16058: waveform_sig_loopback =7277;
16059: waveform_sig_loopback =6285;
16060: waveform_sig_loopback =8277;
16061: waveform_sig_loopback =6939;
16062: waveform_sig_loopback =6160;
16063: waveform_sig_loopback =8349;
16064: waveform_sig_loopback =6757;
16065: waveform_sig_loopback =6822;
16066: waveform_sig_loopback =7169;
16067: waveform_sig_loopback =7918;
16068: waveform_sig_loopback =6416;
16069: waveform_sig_loopback =6500;
16070: waveform_sig_loopback =8592;
16071: waveform_sig_loopback =6644;
16072: waveform_sig_loopback =5735;
16073: waveform_sig_loopback =8327;
16074: waveform_sig_loopback =7759;
16075: waveform_sig_loopback =5492;
16076: waveform_sig_loopback =7193;
16077: waveform_sig_loopback =8655;
16078: waveform_sig_loopback =5488;
16079: waveform_sig_loopback =8719;
16080: waveform_sig_loopback =6118;
16081: waveform_sig_loopback =4370;
16082: waveform_sig_loopback =10134;
16083: waveform_sig_loopback =6837;
16084: waveform_sig_loopback =6382;
16085: waveform_sig_loopback =5960;
16086: waveform_sig_loopback =6943;
16087: waveform_sig_loopback =9033;
16088: waveform_sig_loopback =6002;
16089: waveform_sig_loopback =5883;
16090: waveform_sig_loopback =8046;
16091: waveform_sig_loopback =6049;
16092: waveform_sig_loopback =7823;
16093: waveform_sig_loopback =5995;
16094: waveform_sig_loopback =6607;
16095: waveform_sig_loopback =8207;
16096: waveform_sig_loopback =5503;
16097: waveform_sig_loopback =7242;
16098: waveform_sig_loopback =6898;
16099: waveform_sig_loopback =6649;
16100: waveform_sig_loopback =6240;
16101: waveform_sig_loopback =7587;
16102: waveform_sig_loopback =6445;
16103: waveform_sig_loopback =5952;
16104: waveform_sig_loopback =7558;
16105: waveform_sig_loopback =6509;
16106: waveform_sig_loopback =6251;
16107: waveform_sig_loopback =6531;
16108: waveform_sig_loopback =7645;
16109: waveform_sig_loopback =5663;
16110: waveform_sig_loopback =6050;
16111: waveform_sig_loopback =8223;
16112: waveform_sig_loopback =5736;
16113: waveform_sig_loopback =5326;
16114: waveform_sig_loopback =7933;
16115: waveform_sig_loopback =6785;
16116: waveform_sig_loopback =5107;
16117: waveform_sig_loopback =6587;
16118: waveform_sig_loopback =7754;
16119: waveform_sig_loopback =5156;
16120: waveform_sig_loopback =7943;
16121: waveform_sig_loopback =5188;
16122: waveform_sig_loopback =4101;
16123: waveform_sig_loopback =9136;
16124: waveform_sig_loopback =6327;
16125: waveform_sig_loopback =5553;
16126: waveform_sig_loopback =4990;
16127: waveform_sig_loopback =6648;
16128: waveform_sig_loopback =7884;
16129: waveform_sig_loopback =5207;
16130: waveform_sig_loopback =5349;
16131: waveform_sig_loopback =6837;
16132: waveform_sig_loopback =5371;
16133: waveform_sig_loopback =7123;
16134: waveform_sig_loopback =4951;
16135: waveform_sig_loopback =6026;
16136: waveform_sig_loopback =6926;
16137: waveform_sig_loopback =4762;
16138: waveform_sig_loopback =6669;
16139: waveform_sig_loopback =5627;
16140: waveform_sig_loopback =5757;
16141: waveform_sig_loopback =5538;
16142: waveform_sig_loopback =6583;
16143: waveform_sig_loopback =5517;
16144: waveform_sig_loopback =4925;
16145: waveform_sig_loopback =6467;
16146: waveform_sig_loopback =5884;
16147: waveform_sig_loopback =4834;
16148: waveform_sig_loopback =5663;
16149: waveform_sig_loopback =6793;
16150: waveform_sig_loopback =4199;
16151: waveform_sig_loopback =5390;
16152: waveform_sig_loopback =6939;
16153: waveform_sig_loopback =4531;
16154: waveform_sig_loopback =4626;
16155: waveform_sig_loopback =6517;
16156: waveform_sig_loopback =5754;
16157: waveform_sig_loopback =4137;
16158: waveform_sig_loopback =5303;
16159: waveform_sig_loopback =6727;
16160: waveform_sig_loopback =3930;
16161: waveform_sig_loopback =6825;
16162: waveform_sig_loopback =4001;
16163: waveform_sig_loopback =2949;
16164: waveform_sig_loopback =8004;
16165: waveform_sig_loopback =5249;
16166: waveform_sig_loopback =4092;
16167: waveform_sig_loopback =3921;
16168: waveform_sig_loopback =5681;
16169: waveform_sig_loopback =6366;
16170: waveform_sig_loopback =4184;
16171: waveform_sig_loopback =4063;
16172: waveform_sig_loopback =5571;
16173: waveform_sig_loopback =4600;
16174: waveform_sig_loopback =5326;
16175: waveform_sig_loopback =3806;
16176: waveform_sig_loopback =5136;
16177: waveform_sig_loopback =5410;
16178: waveform_sig_loopback =3645;
16179: waveform_sig_loopback =5171;
16180: waveform_sig_loopback =4330;
16181: waveform_sig_loopback =4853;
16182: waveform_sig_loopback =3813;
16183: waveform_sig_loopback =5281;
16184: waveform_sig_loopback =4391;
16185: waveform_sig_loopback =3379;
16186: waveform_sig_loopback =5388;
16187: waveform_sig_loopback =4338;
16188: waveform_sig_loopback =3359;
16189: waveform_sig_loopback =4779;
16190: waveform_sig_loopback =4998;
16191: waveform_sig_loopback =2884;
16192: waveform_sig_loopback =4371;
16193: waveform_sig_loopback =5230;
16194: waveform_sig_loopback =3238;
16195: waveform_sig_loopback =3234;
16196: waveform_sig_loopback =5042;
16197: waveform_sig_loopback =4512;
16198: waveform_sig_loopback =2393;
16199: waveform_sig_loopback =4016;
16200: waveform_sig_loopback =5451;
16201: waveform_sig_loopback =2233;
16202: waveform_sig_loopback =5540;
16203: waveform_sig_loopback =2290;
16204: waveform_sig_loopback =1572;
16205: waveform_sig_loopback =6756;
16206: waveform_sig_loopback =3543;
16207: waveform_sig_loopback =2484;
16208: waveform_sig_loopback =2683;
16209: waveform_sig_loopback =4014;
16210: waveform_sig_loopback =4872;
16211: waveform_sig_loopback =2835;
16212: waveform_sig_loopback =2219;
16213: waveform_sig_loopback =4171;
16214: waveform_sig_loopback =3001;
16215: waveform_sig_loopback =3686;
16216: waveform_sig_loopback =2587;
16217: waveform_sig_loopback =3096;
16218: waveform_sig_loopback =3816;
16219: waveform_sig_loopback =2368;
16220: waveform_sig_loopback =3216;
16221: waveform_sig_loopback =3107;
16222: waveform_sig_loopback =2975;
16223: waveform_sig_loopback =2092;
16224: waveform_sig_loopback =4113;
16225: waveform_sig_loopback =2250;
16226: waveform_sig_loopback =2070;
16227: waveform_sig_loopback =3780;
16228: waveform_sig_loopback =2369;
16229: waveform_sig_loopback =1964;
16230: waveform_sig_loopback =3026;
16231: waveform_sig_loopback =3230;
16232: waveform_sig_loopback =1250;
16233: waveform_sig_loopback =2613;
16234: waveform_sig_loopback =3484;
16235: waveform_sig_loopback =1641;
16236: waveform_sig_loopback =1442;
16237: waveform_sig_loopback =3384;
16238: waveform_sig_loopback =2832;
16239: waveform_sig_loopback =455;
16240: waveform_sig_loopback =2671;
16241: waveform_sig_loopback =3573;
16242: waveform_sig_loopback =281;
16243: waveform_sig_loopback =4280;
16244: waveform_sig_loopback =14;
16245: waveform_sig_loopback =95;
16246: waveform_sig_loopback =5302;
16247: waveform_sig_loopback =1156;
16248: waveform_sig_loopback =1020;
16249: waveform_sig_loopback =976;
16250: waveform_sig_loopback =2069;
16251: waveform_sig_loopback =3528;
16252: waveform_sig_loopback =465;
16253: waveform_sig_loopback =794;
16254: waveform_sig_loopback =2664;
16255: waveform_sig_loopback =633;
16256: waveform_sig_loopback =2291;
16257: waveform_sig_loopback =482;
16258: waveform_sig_loopback =1430;
16259: waveform_sig_loopback =2308;
16260: waveform_sig_loopback =49;
16261: waveform_sig_loopback =1662;
16262: waveform_sig_loopback =1294;
16263: waveform_sig_loopback =972;
16264: waveform_sig_loopback =512;
16265: waveform_sig_loopback =2125;
16266: waveform_sig_loopback =421;
16267: waveform_sig_loopback =313;
16268: waveform_sig_loopback =1847;
16269: waveform_sig_loopback =605;
16270: waveform_sig_loopback =227;
16271: waveform_sig_loopback =1186;
16272: waveform_sig_loopback =1237;
16273: waveform_sig_loopback =-324;
16274: waveform_sig_loopback =646;
16275: waveform_sig_loopback =1662;
16276: waveform_sig_loopback =-187;
16277: waveform_sig_loopback =-631;
16278: waveform_sig_loopback =1963;
16279: waveform_sig_loopback =578;
16280: waveform_sig_loopback =-1398;
16281: waveform_sig_loopback =1235;
16282: waveform_sig_loopback =1058;
16283: waveform_sig_loopback =-1152;
16284: waveform_sig_loopback =2381;
16285: waveform_sig_loopback =-2328;
16286: waveform_sig_loopback =-1074;
16287: waveform_sig_loopback =2887;
16288: waveform_sig_loopback =-537;
16289: waveform_sig_loopback =-648;
16290: waveform_sig_loopback =-1396;
16291: waveform_sig_loopback =657;
16292: waveform_sig_loopback =1429;
16293: waveform_sig_loopback =-1642;
16294: waveform_sig_loopback =-727;
16295: waveform_sig_loopback =389;
16296: waveform_sig_loopback =-950;
16297: waveform_sig_loopback =469;
16298: waveform_sig_loopback =-1829;
16299: waveform_sig_loopback =26;
16300: waveform_sig_loopback =170;
16301: waveform_sig_loopback =-1822;
16302: waveform_sig_loopback =-123;
16303: waveform_sig_loopback =-842;
16304: waveform_sig_loopback =-724;
16305: waveform_sig_loopback =-1457;
16306: waveform_sig_loopback =252;
16307: waveform_sig_loopback =-1635;
16308: waveform_sig_loopback =-1370;
16309: waveform_sig_loopback =-130;
16310: waveform_sig_loopback =-1402;
16311: waveform_sig_loopback =-1499;
16312: waveform_sig_loopback =-937;
16313: waveform_sig_loopback =-365;
16314: waveform_sig_loopback =-2449;
16315: waveform_sig_loopback =-1308;
16316: waveform_sig_loopback =160;
16317: waveform_sig_loopback =-2592;
16318: waveform_sig_loopback =-2108;
16319: waveform_sig_loopback =67;
16320: waveform_sig_loopback =-1707;
16321: waveform_sig_loopback =-2780;
16322: waveform_sig_loopback =-980;
16323: waveform_sig_loopback =-785;
16324: waveform_sig_loopback =-2785;
16325: waveform_sig_loopback =72;
16326: waveform_sig_loopback =-4020;
16327: waveform_sig_loopback =-2901;
16328: waveform_sig_loopback =896;
16329: waveform_sig_loopback =-2183;
16330: waveform_sig_loopback =-2924;
16331: waveform_sig_loopback =-3048;
16332: waveform_sig_loopback =-1090;
16333: waveform_sig_loopback =-711;
16334: waveform_sig_loopback =-3380;
16335: waveform_sig_loopback =-2628;
16336: waveform_sig_loopback =-1543;
16337: waveform_sig_loopback =-2701;
16338: waveform_sig_loopback =-1528;
16339: waveform_sig_loopback =-3691;
16340: waveform_sig_loopback =-1659;
16341: waveform_sig_loopback =-1878;
16342: waveform_sig_loopback =-3596;
16343: waveform_sig_loopback =-1849;
16344: waveform_sig_loopback =-2746;
16345: waveform_sig_loopback =-2624;
16346: waveform_sig_loopback =-3114;
16347: waveform_sig_loopback =-1800;
16348: waveform_sig_loopback =-3313;
16349: waveform_sig_loopback =-3172;
16350: waveform_sig_loopback =-2151;
16351: waveform_sig_loopback =-2827;
16352: waveform_sig_loopback =-3765;
16353: waveform_sig_loopback =-2419;
16354: waveform_sig_loopback =-2188;
16355: waveform_sig_loopback =-4648;
16356: waveform_sig_loopback =-2467;
16357: waveform_sig_loopback =-2146;
16358: waveform_sig_loopback =-4336;
16359: waveform_sig_loopback =-3595;
16360: waveform_sig_loopback =-2136;
16361: waveform_sig_loopback =-3172;
16362: waveform_sig_loopback =-4772;
16363: waveform_sig_loopback =-2722;
16364: waveform_sig_loopback =-2410;
16365: waveform_sig_loopback =-4807;
16366: waveform_sig_loopback =-1434;
16367: waveform_sig_loopback =-5993;
16368: waveform_sig_loopback =-4531;
16369: waveform_sig_loopback =-695;
16370: waveform_sig_loopback =-4174;
16371: waveform_sig_loopback =-4662;
16372: waveform_sig_loopback =-4573;
16373: waveform_sig_loopback =-2815;
16374: waveform_sig_loopback =-2526;
16375: waveform_sig_loopback =-5056;
16376: waveform_sig_loopback =-4215;
16377: waveform_sig_loopback =-3330;
16378: waveform_sig_loopback =-4246;
16379: waveform_sig_loopback =-3418;
16380: waveform_sig_loopback =-5208;
16381: waveform_sig_loopback =-3206;
16382: waveform_sig_loopback =-3903;
16383: waveform_sig_loopback =-4935;
16384: waveform_sig_loopback =-3672;
16385: waveform_sig_loopback =-4445;
16386: waveform_sig_loopback =-4041;
16387: waveform_sig_loopback =-5075;
16388: waveform_sig_loopback =-3168;
16389: waveform_sig_loopback =-5005;
16390: waveform_sig_loopback =-4997;
16391: waveform_sig_loopback =-3455;
16392: waveform_sig_loopback =-4788;
16393: waveform_sig_loopback =-5257;
16394: waveform_sig_loopback =-3802;
16395: waveform_sig_loopback =-4260;
16396: waveform_sig_loopback =-5916;
16397: waveform_sig_loopback =-4065;
16398: waveform_sig_loopback =-3875;
16399: waveform_sig_loopback =-5777;
16400: waveform_sig_loopback =-5238;
16401: waveform_sig_loopback =-3593;
16402: waveform_sig_loopback =-4768;
16403: waveform_sig_loopback =-6442;
16404: waveform_sig_loopback =-4044;
16405: waveform_sig_loopback =-3993;
16406: waveform_sig_loopback =-6410;
16407: waveform_sig_loopback =-2807;
16408: waveform_sig_loopback =-7725;
16409: waveform_sig_loopback =-5857;
16410: waveform_sig_loopback =-2111;
16411: waveform_sig_loopback =-5902;
16412: waveform_sig_loopback =-6144;
16413: waveform_sig_loopback =-5845;
16414: waveform_sig_loopback =-4437;
16415: waveform_sig_loopback =-3935;
16416: waveform_sig_loopback =-6560;
16417: waveform_sig_loopback =-5722;
16418: waveform_sig_loopback =-4619;
16419: waveform_sig_loopback =-5733;
16420: waveform_sig_loopback =-4917;
16421: waveform_sig_loopback =-6425;
16422: waveform_sig_loopback =-4811;
16423: waveform_sig_loopback =-5209;
16424: waveform_sig_loopback =-6184;
16425: waveform_sig_loopback =-5291;
16426: waveform_sig_loopback =-5561;
16427: waveform_sig_loopback =-5585;
16428: waveform_sig_loopback =-6473;
16429: waveform_sig_loopback =-4157;
16430: waveform_sig_loopback =-6794;
16431: waveform_sig_loopback =-6110;
16432: waveform_sig_loopback =-4694;
16433: waveform_sig_loopback =-6372;
16434: waveform_sig_loopback =-6235;
16435: waveform_sig_loopback =-5227;
16436: waveform_sig_loopback =-5600;
16437: waveform_sig_loopback =-7017;
16438: waveform_sig_loopback =-5443;
16439: waveform_sig_loopback =-5056;
16440: waveform_sig_loopback =-7073;
16441: waveform_sig_loopback =-6490;
16442: waveform_sig_loopback =-4640;
16443: waveform_sig_loopback =-6069;
16444: waveform_sig_loopback =-7762;
16445: waveform_sig_loopback =-4904;
16446: waveform_sig_loopback =-5416;
16447: waveform_sig_loopback =-7518;
16448: waveform_sig_loopback =-3792;
16449: waveform_sig_loopback =-9263;
16450: waveform_sig_loopback =-6536;
16451: waveform_sig_loopback =-3261;
16452: waveform_sig_loopback =-7316;
16453: waveform_sig_loopback =-6960;
16454: waveform_sig_loopback =-7029;
16455: waveform_sig_loopback =-5572;
16456: waveform_sig_loopback =-4812;
16457: waveform_sig_loopback =-8026;
16458: waveform_sig_loopback =-6509;
16459: waveform_sig_loopback =-5634;
16460: waveform_sig_loopback =-7064;
16461: waveform_sig_loopback =-5682;
16462: waveform_sig_loopback =-7649;
16463: waveform_sig_loopback =-5742;
16464: waveform_sig_loopback =-6162;
16465: waveform_sig_loopback =-7424;
16466: waveform_sig_loopback =-6154;
16467: waveform_sig_loopback =-6459;
16468: waveform_sig_loopback =-6782;
16469: waveform_sig_loopback =-7200;
16470: waveform_sig_loopback =-5198;
16471: waveform_sig_loopback =-7894;
16472: waveform_sig_loopback =-6687;
16473: waveform_sig_loopback =-5793;
16474: waveform_sig_loopback =-7362;
16475: waveform_sig_loopback =-6917;
16476: waveform_sig_loopback =-6361;
16477: waveform_sig_loopback =-6344;
16478: waveform_sig_loopback =-7846;
16479: waveform_sig_loopback =-6463;
16480: waveform_sig_loopback =-5799;
16481: waveform_sig_loopback =-8122;
16482: waveform_sig_loopback =-7087;
16483: waveform_sig_loopback =-5340;
16484: waveform_sig_loopback =-7408;
16485: waveform_sig_loopback =-8289;
16486: waveform_sig_loopback =-5449;
16487: waveform_sig_loopback =-6507;
16488: waveform_sig_loopback =-8096;
16489: waveform_sig_loopback =-4749;
16490: waveform_sig_loopback =-10032;
16491: waveform_sig_loopback =-6865;
16492: waveform_sig_loopback =-4420;
16493: waveform_sig_loopback =-8027;
16494: waveform_sig_loopback =-7471;
16495: waveform_sig_loopback =-7992;
16496: waveform_sig_loopback =-6014;
16497: waveform_sig_loopback =-5587;
16498: waveform_sig_loopback =-8851;
16499: waveform_sig_loopback =-6848;
16500: waveform_sig_loopback =-6651;
16501: waveform_sig_loopback =-7521;
16502: waveform_sig_loopback =-6128;
16503: waveform_sig_loopback =-8595;
16504: waveform_sig_loopback =-6110;
16505: waveform_sig_loopback =-6785;
16506: waveform_sig_loopback =-8111;
16507: waveform_sig_loopback =-6527;
16508: waveform_sig_loopback =-7185;
16509: waveform_sig_loopback =-7364;
16510: waveform_sig_loopback =-7367;
16511: waveform_sig_loopback =-6118;
16512: waveform_sig_loopback =-8269;
16513: waveform_sig_loopback =-6948;
16514: waveform_sig_loopback =-6597;
16515: waveform_sig_loopback =-7520;
16516: waveform_sig_loopback =-7628;
16517: waveform_sig_loopback =-6628;
16518: waveform_sig_loopback =-6716;
16519: waveform_sig_loopback =-8561;
16520: waveform_sig_loopback =-6626;
16521: waveform_sig_loopback =-6082;
16522: waveform_sig_loopback =-8681;
16523: waveform_sig_loopback =-7391;
16524: waveform_sig_loopback =-5726;
16525: waveform_sig_loopback =-7685;
16526: waveform_sig_loopback =-8486;
16527: waveform_sig_loopback =-5949;
16528: waveform_sig_loopback =-6981;
16529: waveform_sig_loopback =-7978;
16530: waveform_sig_loopback =-5223;
16531: waveform_sig_loopback =-10647;
16532: waveform_sig_loopback =-6672;
16533: waveform_sig_loopback =-4943;
16534: waveform_sig_loopback =-8072;
16535: waveform_sig_loopback =-7864;
16536: waveform_sig_loopback =-8294;
16537: waveform_sig_loopback =-5724;
16538: waveform_sig_loopback =-6232;
16539: waveform_sig_loopback =-8961;
16540: waveform_sig_loopback =-6752;
16541: waveform_sig_loopback =-7098;
16542: waveform_sig_loopback =-7324;
16543: waveform_sig_loopback =-6587;
16544: waveform_sig_loopback =-8641;
16545: waveform_sig_loopback =-5854;
16546: waveform_sig_loopback =-7356;
16547: waveform_sig_loopback =-7909;
16548: waveform_sig_loopback =-6548;
16549: waveform_sig_loopback =-7368;
16550: waveform_sig_loopback =-7289;
16551: waveform_sig_loopback =-7466;
16552: waveform_sig_loopback =-6139;
16553: waveform_sig_loopback =-8184;
16554: waveform_sig_loopback =-7060;
16555: waveform_sig_loopback =-6562;
16556: waveform_sig_loopback =-7417;
16557: waveform_sig_loopback =-7709;
16558: waveform_sig_loopback =-6433;
16559: waveform_sig_loopback =-6766;
16560: waveform_sig_loopback =-8532;
16561: waveform_sig_loopback =-6240;
16562: waveform_sig_loopback =-6281;
16563: waveform_sig_loopback =-8591;
16564: waveform_sig_loopback =-6995;
16565: waveform_sig_loopback =-5722;
16566: waveform_sig_loopback =-7641;
16567: waveform_sig_loopback =-8168;
16568: waveform_sig_loopback =-5834;
16569: waveform_sig_loopback =-6852;
16570: waveform_sig_loopback =-7668;
16571: waveform_sig_loopback =-5297;
16572: waveform_sig_loopback =-10234;
16573: waveform_sig_loopback =-6395;
16574: waveform_sig_loopback =-4848;
16575: waveform_sig_loopback =-7574;
16576: waveform_sig_loopback =-8009;
16577: waveform_sig_loopback =-7655;
16578: waveform_sig_loopback =-5429;
16579: waveform_sig_loopback =-6242;
16580: waveform_sig_loopback =-8275;
16581: waveform_sig_loopback =-6686;
16582: waveform_sig_loopback =-6662;
16583: waveform_sig_loopback =-6804;
16584: waveform_sig_loopback =-6594;
16585: waveform_sig_loopback =-7941;
16586: waveform_sig_loopback =-5559;
16587: waveform_sig_loopback =-7122;
16588: waveform_sig_loopback =-7218;
16589: waveform_sig_loopback =-6375;
16590: waveform_sig_loopback =-6841;
16591: waveform_sig_loopback =-6827;
16592: waveform_sig_loopback =-7034;
16593: waveform_sig_loopback =-5693;
16594: waveform_sig_loopback =-7723;
16595: waveform_sig_loopback =-6583;
16596: waveform_sig_loopback =-6040;
16597: waveform_sig_loopback =-6874;
16598: waveform_sig_loopback =-7339;
16599: waveform_sig_loopback =-5625;
16600: waveform_sig_loopback =-6464;
16601: waveform_sig_loopback =-7998;
16602: waveform_sig_loopback =-5331;
16603: waveform_sig_loopback =-6154;
16604: waveform_sig_loopback =-7771;
16605: waveform_sig_loopback =-6279;
16606: waveform_sig_loopback =-5450;
16607: waveform_sig_loopback =-6703;
16608: waveform_sig_loopback =-7786;
16609: waveform_sig_loopback =-5049;
16610: waveform_sig_loopback =-6120;
16611: waveform_sig_loopback =-7184;
16612: waveform_sig_loopback =-4380;
16613: waveform_sig_loopback =-9732;
16614: waveform_sig_loopback =-5553;
16615: waveform_sig_loopback =-3911;
16616: waveform_sig_loopback =-7218;
16617: waveform_sig_loopback =-7174;
16618: waveform_sig_loopback =-6658;
16619: waveform_sig_loopback =-4957;
16620: waveform_sig_loopback =-5308;
16621: waveform_sig_loopback =-7601;
16622: waveform_sig_loopback =-5906;
16623: waveform_sig_loopback =-5747;
16624: waveform_sig_loopback =-6130;
16625: waveform_sig_loopback =-5738;
16626: waveform_sig_loopback =-6978;
16627: waveform_sig_loopback =-4825;
16628: waveform_sig_loopback =-6269;
16629: waveform_sig_loopback =-6250;
16630: waveform_sig_loopback =-5615;
16631: waveform_sig_loopback =-5866;
16632: waveform_sig_loopback =-5928;
16633: waveform_sig_loopback =-6248;
16634: waveform_sig_loopback =-4561;
16635: waveform_sig_loopback =-6921;
16636: waveform_sig_loopback =-5686;
16637: waveform_sig_loopback =-4774;
16638: waveform_sig_loopback =-6346;
16639: waveform_sig_loopback =-6048;
16640: waveform_sig_loopback =-4566;
16641: waveform_sig_loopback =-5906;
16642: waveform_sig_loopback =-6409;
16643: waveform_sig_loopback =-4650;
16644: waveform_sig_loopback =-5073;
16645: waveform_sig_loopback =-6566;
16646: waveform_sig_loopback =-5527;
16647: waveform_sig_loopback =-4005;
16648: waveform_sig_loopback =-5946;
16649: waveform_sig_loopback =-6703;
16650: waveform_sig_loopback =-3683;
16651: waveform_sig_loopback =-5409;
16652: waveform_sig_loopback =-5837;
16653: waveform_sig_loopback =-3362;
16654: waveform_sig_loopback =-8785;
16655: waveform_sig_loopback =-4154;
16656: waveform_sig_loopback =-2869;
16657: waveform_sig_loopback =-6209;
16658: waveform_sig_loopback =-5891;
16659: waveform_sig_loopback =-5461;
16660: waveform_sig_loopback =-3819;
16661: waveform_sig_loopback =-3959;
16662: waveform_sig_loopback =-6629;
16663: waveform_sig_loopback =-4627;
16664: waveform_sig_loopback =-4393;
16665: waveform_sig_loopback =-5083;
16666: waveform_sig_loopback =-4385;
16667: waveform_sig_loopback =-5722;
16668: waveform_sig_loopback =-3737;
16669: waveform_sig_loopback =-4780;
16670: waveform_sig_loopback =-5083;
16671: waveform_sig_loopback =-4404;
16672: waveform_sig_loopback =-4283;
16673: waveform_sig_loopback =-4999;
16674: waveform_sig_loopback =-4605;
16675: waveform_sig_loopback =-3257;
16676: waveform_sig_loopback =-5904;
16677: waveform_sig_loopback =-3833;
16678: waveform_sig_loopback =-3717;
16679: waveform_sig_loopback =-5015;
16680: waveform_sig_loopback =-4411;
16681: waveform_sig_loopback =-3465;
16682: waveform_sig_loopback =-4320;
16683: waveform_sig_loopback =-5038;
16684: waveform_sig_loopback =-3373;
16685: waveform_sig_loopback =-3470;
16686: waveform_sig_loopback =-5328;
16687: waveform_sig_loopback =-3997;
16688: waveform_sig_loopback =-2452;
16689: waveform_sig_loopback =-4742;
16690: waveform_sig_loopback =-5043;
16691: waveform_sig_loopback =-2081;
16692: waveform_sig_loopback =-4288;
16693: waveform_sig_loopback =-3986;
16694: waveform_sig_loopback =-2004;
16695: waveform_sig_loopback =-7518;
16696: waveform_sig_loopback =-2131;
16697: waveform_sig_loopback =-1664;
16698: waveform_sig_loopback =-4766;
16699: waveform_sig_loopback =-4144;
16700: waveform_sig_loopback =-4199;
16701: waveform_sig_loopback =-2026;
16702: waveform_sig_loopback =-2426;
16703: waveform_sig_loopback =-5419;
16704: waveform_sig_loopback =-2555;
16705: waveform_sig_loopback =-3128;
16706: waveform_sig_loopback =-3490;
16707: waveform_sig_loopback =-2565;
16708: waveform_sig_loopback =-4532;
16709: waveform_sig_loopback =-1731;
16710: waveform_sig_loopback =-3293;
16711: waveform_sig_loopback =-3715;
16712: waveform_sig_loopback =-2413;
16713: waveform_sig_loopback =-2963;
16714: waveform_sig_loopback =-3352;
16715: waveform_sig_loopback =-2701;
16716: waveform_sig_loopback =-2032;
16717: waveform_sig_loopback =-3979;
16718: waveform_sig_loopback =-2208;
16719: waveform_sig_loopback =-2282;
16720: waveform_sig_loopback =-3113;
16721: waveform_sig_loopback =-2878;
16722: waveform_sig_loopback =-1731;
16723: waveform_sig_loopback =-2699;
16724: waveform_sig_loopback =-3394;
16725: waveform_sig_loopback =-1573;
16726: waveform_sig_loopback =-1813;
16727: waveform_sig_loopback =-3736;
16728: waveform_sig_loopback =-2192;
16729: waveform_sig_loopback =-607;
16730: waveform_sig_loopback =-3386;
16731: waveform_sig_loopback =-3046;
16732: waveform_sig_loopback =-321;
16733: waveform_sig_loopback =-2915;
16734: waveform_sig_loopback =-1683;
16735: waveform_sig_loopback =-914;
16736: waveform_sig_loopback =-5579;
16737: waveform_sig_loopback =35;
16738: waveform_sig_loopback =-594;
16739: waveform_sig_loopback =-2449;
16740: waveform_sig_loopback =-2682;
16741: waveform_sig_loopback =-2419;
16742: waveform_sig_loopback =196;
16743: waveform_sig_loopback =-1305;
16744: waveform_sig_loopback =-3184;
16745: waveform_sig_loopback =-755;
16746: waveform_sig_loopback =-1715;
16747: waveform_sig_loopback =-1186;
16748: waveform_sig_loopback =-1205;
16749: waveform_sig_loopback =-2571;
16750: waveform_sig_loopback =298;
16751: waveform_sig_loopback =-1925;
16752: waveform_sig_loopback =-1530;
16753: waveform_sig_loopback =-762;
16754: waveform_sig_loopback =-1171;
16755: waveform_sig_loopback =-1441;
16756: waveform_sig_loopback =-908;
16757: waveform_sig_loopback =-252;
16758: waveform_sig_loopback =-2158;
16759: waveform_sig_loopback =-219;
16760: waveform_sig_loopback =-664;
16761: waveform_sig_loopback =-1071;
16762: waveform_sig_loopback =-1174;
16763: waveform_sig_loopback =150;
16764: waveform_sig_loopback =-619;
16765: waveform_sig_loopback =-1966;
16766: waveform_sig_loopback =740;
16767: waveform_sig_loopback =-195;
16768: waveform_sig_loopback =-2066;
16769: waveform_sig_loopback =198;
16770: waveform_sig_loopback =695;
16771: waveform_sig_loopback =-1316;
16772: waveform_sig_loopback =-965;
16773: waveform_sig_loopback =1185;
16774: waveform_sig_loopback =-664;
16775: waveform_sig_loopback =87;
16776: waveform_sig_loopback =787;
16777: waveform_sig_loopback =-3366;
16778: waveform_sig_loopback =1761;
16779: waveform_sig_loopback =1462;
16780: waveform_sig_loopback =-542;
16781: waveform_sig_loopback =-1147;
16782: waveform_sig_loopback =-6;
16783: waveform_sig_loopback =1866;
16784: waveform_sig_loopback =531;
16785: waveform_sig_loopback =-1161;
16786: waveform_sig_loopback =964;
16787: waveform_sig_loopback =342;
16788: waveform_sig_loopback =781;
16789: waveform_sig_loopback =466;
16790: waveform_sig_loopback =-466;
16791: waveform_sig_loopback =2166;
16792: waveform_sig_loopback =-183;
16793: waveform_sig_loopback =563;
16794: waveform_sig_loopback =1107;
16795: waveform_sig_loopback =677;
16796: waveform_sig_loopback =649;
16797: waveform_sig_loopback =951;
16798: waveform_sig_loopback =1574;
16799: waveform_sig_loopback =-38;
16800: waveform_sig_loopback =1437;
16801: waveform_sig_loopback =1556;
16802: waveform_sig_loopback =745;
16803: waveform_sig_loopback =473;
16804: waveform_sig_loopback =2560;
16805: waveform_sig_loopback =694;
16806: waveform_sig_loopback =204;
16807: waveform_sig_loopback =2908;
16808: waveform_sig_loopback =1230;
16809: waveform_sig_loopback =303;
16810: waveform_sig_loopback =1961;
16811: waveform_sig_loopback =2486;
16812: waveform_sig_loopback =866;
16813: waveform_sig_loopback =603;
16814: waveform_sig_loopback =3362;
16815: waveform_sig_loopback =1149;
16816: waveform_sig_loopback =1888;
16817: waveform_sig_loopback =2870;
16818: waveform_sig_loopback =-1733;
16819: waveform_sig_loopback =3830;
16820: waveform_sig_loopback =3439;
16821: waveform_sig_loopback =884;
16822: waveform_sig_loopback =1059;
16823: waveform_sig_loopback =1906;
16824: waveform_sig_loopback =3596;
16825: waveform_sig_loopback =2420;
16826: waveform_sig_loopback =602;
16827: waveform_sig_loopback =2966;
16828: waveform_sig_loopback =2106;
16829: waveform_sig_loopback =2651;
16830: waveform_sig_loopback =1998;
16831: waveform_sig_loopback =1716;
16832: waveform_sig_loopback =3941;
16833: waveform_sig_loopback =1487;
16834: waveform_sig_loopback =2507;
16835: waveform_sig_loopback =2619;
16836: waveform_sig_loopback =2922;
16837: waveform_sig_loopback =2329;
16838: waveform_sig_loopback =2433;
16839: waveform_sig_loopback =3806;
16840: waveform_sig_loopback =1509;
16841: waveform_sig_loopback =3292;
16842: waveform_sig_loopback =3425;
16843: waveform_sig_loopback =2030;
16844: waveform_sig_loopback =3044;
16845: waveform_sig_loopback =3951;
16846: waveform_sig_loopback =2270;
16847: waveform_sig_loopback =2498;
16848: waveform_sig_loopback =4233;
16849: waveform_sig_loopback =3216;
16850: waveform_sig_loopback =1873;
16851: waveform_sig_loopback =3770;
16852: waveform_sig_loopback =4497;
16853: waveform_sig_loopback =2269;
16854: waveform_sig_loopback =2446;
16855: waveform_sig_loopback =5281;
16856: waveform_sig_loopback =2668;
16857: waveform_sig_loopback =3748;
16858: waveform_sig_loopback =4474;
16859: waveform_sig_loopback =-44;
16860: waveform_sig_loopback =5849;
16861: waveform_sig_loopback =4967;
16862: waveform_sig_loopback =2445;
16863: waveform_sig_loopback =2959;
16864: waveform_sig_loopback =3552;
16865: waveform_sig_loopback =5229;
16866: waveform_sig_loopback =4199;
16867: waveform_sig_loopback =2226;
16868: waveform_sig_loopback =4709;
16869: waveform_sig_loopback =3889;
16870: waveform_sig_loopback =4136;
16871: waveform_sig_loopback =3981;
16872: waveform_sig_loopback =3336;
16873: waveform_sig_loopback =5291;
16874: waveform_sig_loopback =3484;
16875: waveform_sig_loopback =4124;
16876: waveform_sig_loopback =4263;
16877: waveform_sig_loopback =4583;
16878: waveform_sig_loopback =3557;
16879: waveform_sig_loopback =4671;
16880: waveform_sig_loopback =5191;
16881: waveform_sig_loopback =2803;
16882: waveform_sig_loopback =5429;
16883: waveform_sig_loopback =4716;
16884: waveform_sig_loopback =3771;
16885: waveform_sig_loopback =4567;
16886: waveform_sig_loopback =5310;
16887: waveform_sig_loopback =4218;
16888: waveform_sig_loopback =3845;
16889: waveform_sig_loopback =5798;
16890: waveform_sig_loopback =4896;
16891: waveform_sig_loopback =3313;
16892: waveform_sig_loopback =5454;
16893: waveform_sig_loopback =5943;
16894: waveform_sig_loopback =3702;
16895: waveform_sig_loopback =4191;
16896: waveform_sig_loopback =6847;
16897: waveform_sig_loopback =3873;
16898: waveform_sig_loopback =5622;
16899: waveform_sig_loopback =5746;
16900: waveform_sig_loopback =1323;
16901: waveform_sig_loopback =7699;
16902: waveform_sig_loopback =6091;
16903: waveform_sig_loopback =3985;
16904: waveform_sig_loopback =4514;
16905: waveform_sig_loopback =4751;
16906: waveform_sig_loopback =7018;
16907: waveform_sig_loopback =5413;
16908: waveform_sig_loopback =3511;
16909: waveform_sig_loopback =6425;
16910: waveform_sig_loopback =5058;
16911: waveform_sig_loopback =5659;
16912: waveform_sig_loopback =5379;
16913: waveform_sig_loopback =4580;
16914: waveform_sig_loopback =6894;
16915: waveform_sig_loopback =4776;
16916: waveform_sig_loopback =5340;
16917: waveform_sig_loopback =5956;
16918: waveform_sig_loopback =5736;
16919: waveform_sig_loopback =4863;
16920: waveform_sig_loopback =6350;
16921: waveform_sig_loopback =6083;
16922: waveform_sig_loopback =4435;
16923: waveform_sig_loopback =6733;
16924: waveform_sig_loopback =5776;
16925: waveform_sig_loopback =5387;
16926: waveform_sig_loopback =5684;
16927: waveform_sig_loopback =6677;
16928: waveform_sig_loopback =5489;
16929: waveform_sig_loopback =5005;
16930: waveform_sig_loopback =7246;
16931: waveform_sig_loopback =5934;
16932: waveform_sig_loopback =4523;
16933: waveform_sig_loopback =6878;
16934: waveform_sig_loopback =7023;
16935: waveform_sig_loopback =4784;
16936: waveform_sig_loopback =5612;
16937: waveform_sig_loopback =7908;
16938: waveform_sig_loopback =4884;
16939: waveform_sig_loopback =7177;
16940: waveform_sig_loopback =6444;
16941: waveform_sig_loopback =2749;
16942: waveform_sig_loopback =9115;
16943: waveform_sig_loopback =6804;
16944: waveform_sig_loopback =5450;
16945: waveform_sig_loopback =5412;
16946: waveform_sig_loopback =5963;
16947: waveform_sig_loopback =8374;
16948: waveform_sig_loopback =6053;
16949: waveform_sig_loopback =4942;
16950: waveform_sig_loopback =7536;
16951: waveform_sig_loopback =5827;
16952: waveform_sig_loopback =7098;
16953: waveform_sig_loopback =6105;
16954: waveform_sig_loopback =5736;
16955: waveform_sig_loopback =8110;
16956: waveform_sig_loopback =5452;
16957: waveform_sig_loopback =6664;
16958: waveform_sig_loopback =6903;
16959: waveform_sig_loopback =6521;
16960: waveform_sig_loopback =6099;
16961: waveform_sig_loopback =7208;
16962: waveform_sig_loopback =6907;
16963: waveform_sig_loopback =5627;
16964: waveform_sig_loopback =7450;
16965: waveform_sig_loopback =6803;
16966: waveform_sig_loopback =6342;
16967: waveform_sig_loopback =6406;
16968: waveform_sig_loopback =7833;
16969: waveform_sig_loopback =6178;
16970: waveform_sig_loopback =5900;
16971: waveform_sig_loopback =8334;
16972: waveform_sig_loopback =6484;
16973: waveform_sig_loopback =5520;
16974: waveform_sig_loopback =7838;
16975: waveform_sig_loopback =7623;
16976: waveform_sig_loopback =5702;
16977: waveform_sig_loopback =6474;
16978: waveform_sig_loopback =8584;
16979: waveform_sig_loopback =5735;
16980: waveform_sig_loopback =8035;
16981: waveform_sig_loopback =6809;
16982: waveform_sig_loopback =3821;
16983: waveform_sig_loopback =9759;
16984: waveform_sig_loopback =7428;
16985: waveform_sig_loopback =6309;
16986: waveform_sig_loopback =5838;
16987: waveform_sig_loopback =7028;
16988: waveform_sig_loopback =8933;
16989: waveform_sig_loopback =6440;
16990: waveform_sig_loopback =5989;
16991: waveform_sig_loopback =7840;
16992: waveform_sig_loopback =6588;
16993: waveform_sig_loopback =7894;
16994: waveform_sig_loopback =6288;
16995: waveform_sig_loopback =6797;
16996: waveform_sig_loopback =8431;
16997: waveform_sig_loopback =5882;
16998: waveform_sig_loopback =7527;
16999: waveform_sig_loopback =7043;
17000: waveform_sig_loopback =7305;
17001: waveform_sig_loopback =6615;
17002: waveform_sig_loopback =7565;
17003: waveform_sig_loopback =7581;
17004: waveform_sig_loopback =5966;
17005: waveform_sig_loopback =8000;
17006: waveform_sig_loopback =7315;
17007: waveform_sig_loopback =6578;
17008: waveform_sig_loopback =7060;
17009: waveform_sig_loopback =8239;
17010: waveform_sig_loopback =6394;
17011: waveform_sig_loopback =6452;
17012: waveform_sig_loopback =8761;
17013: waveform_sig_loopback =6715;
17014: waveform_sig_loopback =5959;
17015: waveform_sig_loopback =8296;
17016: waveform_sig_loopback =7741;
17017: waveform_sig_loopback =6161;
17018: waveform_sig_loopback =6803;
17019: waveform_sig_loopback =8790;
17020: waveform_sig_loopback =6206;
17021: waveform_sig_loopback =8139;
17022: waveform_sig_loopback =7124;
17023: waveform_sig_loopback =4238;
17024: waveform_sig_loopback =9808;
17025: waveform_sig_loopback =7977;
17026: waveform_sig_loopback =6178;
17027: waveform_sig_loopback =6130;
17028: waveform_sig_loopback =7527;
17029: waveform_sig_loopback =8697;
17030: waveform_sig_loopback =6958;
17031: waveform_sig_loopback =6013;
17032: waveform_sig_loopback =7913;
17033: waveform_sig_loopback =7042;
17034: waveform_sig_loopback =7673;
17035: waveform_sig_loopback =6584;
17036: waveform_sig_loopback =7062;
17037: waveform_sig_loopback =8243;
17038: waveform_sig_loopback =6265;
17039: waveform_sig_loopback =7449;
17040: waveform_sig_loopback =7129;
17041: waveform_sig_loopback =7445;
17042: waveform_sig_loopback =6462;
17043: waveform_sig_loopback =7828;
17044: waveform_sig_loopback =7438;
17045: waveform_sig_loopback =6005;
17046: waveform_sig_loopback =7996;
17047: waveform_sig_loopback =7354;
17048: waveform_sig_loopback =6422;
17049: waveform_sig_loopback =7111;
17050: waveform_sig_loopback =8293;
17051: waveform_sig_loopback =6012;
17052: waveform_sig_loopback =6797;
17053: waveform_sig_loopback =8472;
17054: waveform_sig_loopback =6447;
17055: waveform_sig_loopback =6220;
17056: waveform_sig_loopback =7873;
17057: waveform_sig_loopback =7818;
17058: waveform_sig_loopback =5947;
17059: waveform_sig_loopback =6501;
17060: waveform_sig_loopback =8991;
17061: waveform_sig_loopback =5597;
17062: waveform_sig_loopback =8170;
17063: waveform_sig_loopback =6858;
17064: waveform_sig_loopback =3782;
17065: waveform_sig_loopback =10050;
17066: waveform_sig_loopback =7449;
17067: waveform_sig_loopback =5715;
17068: waveform_sig_loopback =6308;
17069: waveform_sig_loopback =6961;
17070: waveform_sig_loopback =8511;
17071: waveform_sig_loopback =6668;
17072: waveform_sig_loopback =5475;
17073: waveform_sig_loopback =7927;
17074: waveform_sig_loopback =6469;
17075: waveform_sig_loopback =7291;
17076: waveform_sig_loopback =6404;
17077: waveform_sig_loopback =6516;
17078: waveform_sig_loopback =7897;
17079: waveform_sig_loopback =5873;
17080: waveform_sig_loopback =6982;
17081: waveform_sig_loopback =6776;
17082: waveform_sig_loopback =6950;
17083: waveform_sig_loopback =5989;
17084: waveform_sig_loopback =7411;
17085: waveform_sig_loopback =6980;
17086: waveform_sig_loopback =5411;
17087: waveform_sig_loopback =7649;
17088: waveform_sig_loopback =6826;
17089: waveform_sig_loopback =5672;
17090: waveform_sig_loopback =7032;
17091: waveform_sig_loopback =7330;
17092: waveform_sig_loopback =5534;
17093: waveform_sig_loopback =6507;
17094: waveform_sig_loopback =7422;
17095: waveform_sig_loopback =6317;
17096: waveform_sig_loopback =5336;
17097: waveform_sig_loopback =7281;
17098: waveform_sig_loopback =7494;
17099: waveform_sig_loopback =4725;
17100: waveform_sig_loopback =6450;
17101: waveform_sig_loopback =8132;
17102: waveform_sig_loopback =4672;
17103: waveform_sig_loopback =8095;
17104: waveform_sig_loopback =5452;
17105: waveform_sig_loopback =3540;
17106: waveform_sig_loopback =9429;
17107: waveform_sig_loopback =6322;
17108: waveform_sig_loopback =5345;
17109: waveform_sig_loopback =5281;
17110: waveform_sig_loopback =6351;
17111: waveform_sig_loopback =7866;
17112: waveform_sig_loopback =5636;
17113: waveform_sig_loopback =4830;
17114: waveform_sig_loopback =7140;
17115: waveform_sig_loopback =5653;
17116: waveform_sig_loopback =6461;
17117: waveform_sig_loopback =5505;
17118: waveform_sig_loopback =5710;
17119: waveform_sig_loopback =7035;
17120: waveform_sig_loopback =5076;
17121: waveform_sig_loopback =5978;
17122: waveform_sig_loopback =6073;
17123: waveform_sig_loopback =6101;
17124: waveform_sig_loopback =4829;
17125: waveform_sig_loopback =6900;
17126: waveform_sig_loopback =5637;
17127: waveform_sig_loopback =4728;
17128: waveform_sig_loopback =6871;
17129: waveform_sig_loopback =5341;
17130: waveform_sig_loopback =5231;
17131: waveform_sig_loopback =5865;
17132: waveform_sig_loopback =6264;
17133: waveform_sig_loopback =4837;
17134: waveform_sig_loopback =5149;
17135: waveform_sig_loopback =6818;
17136: waveform_sig_loopback =5087;
17137: waveform_sig_loopback =4193;
17138: waveform_sig_loopback =6655;
17139: waveform_sig_loopback =6056;
17140: waveform_sig_loopback =3755;
17141: waveform_sig_loopback =5552;
17142: waveform_sig_loopback =6808;
17143: waveform_sig_loopback =3752;
17144: waveform_sig_loopback =7054;
17145: waveform_sig_loopback =4029;
17146: waveform_sig_loopback =2754;
17147: waveform_sig_loopback =8277;
17148: waveform_sig_loopback =5030;
17149: waveform_sig_loopback =4236;
17150: waveform_sig_loopback =4069;
17151: waveform_sig_loopback =5175;
17152: waveform_sig_loopback =6810;
17153: waveform_sig_loopback =4212;
17154: waveform_sig_loopback =3660;
17155: waveform_sig_loopback =6104;
17156: waveform_sig_loopback =4108;
17157: waveform_sig_loopback =5567;
17158: waveform_sig_loopback =4070;
17159: waveform_sig_loopback =4376;
17160: waveform_sig_loopback =6103;
17161: waveform_sig_loopback =3416;
17162: waveform_sig_loopback =4891;
17163: waveform_sig_loopback =4839;
17164: waveform_sig_loopback =4383;
17165: waveform_sig_loopback =3995;
17166: waveform_sig_loopback =5442;
17167: waveform_sig_loopback =4068;
17168: waveform_sig_loopback =3760;
17169: waveform_sig_loopback =5217;
17170: waveform_sig_loopback =4232;
17171: waveform_sig_loopback =3853;
17172: waveform_sig_loopback =4329;
17173: waveform_sig_loopback =5166;
17174: waveform_sig_loopback =3121;
17175: waveform_sig_loopback =3861;
17176: waveform_sig_loopback =5503;
17177: waveform_sig_loopback =3429;
17178: waveform_sig_loopback =2888;
17179: waveform_sig_loopback =5105;
17180: waveform_sig_loopback =4583;
17181: waveform_sig_loopback =2372;
17182: waveform_sig_loopback =4248;
17183: waveform_sig_loopback =4915;
17184: waveform_sig_loopback =2477;
17185: waveform_sig_loopback =5875;
17186: waveform_sig_loopback =2006;
17187: waveform_sig_loopback =1613;
17188: waveform_sig_loopback =6673;
17189: waveform_sig_loopback =3571;
17190: waveform_sig_loopback =2836;
17191: waveform_sig_loopback =2172;
17192: waveform_sig_loopback =4057;
17193: waveform_sig_loopback =5276;
17194: waveform_sig_loopback =2235;
17195: waveform_sig_loopback =2540;
17196: waveform_sig_loopback =4294;
17197: waveform_sig_loopback =2596;
17198: waveform_sig_loopback =4193;
17199: waveform_sig_loopback =1986;
17200: waveform_sig_loopback =3376;
17201: waveform_sig_loopback =4313;
17202: waveform_sig_loopback =1617;
17203: waveform_sig_loopback =3696;
17204: waveform_sig_loopback =2891;
17205: waveform_sig_loopback =3017;
17206: waveform_sig_loopback =2344;
17207: waveform_sig_loopback =3566;
17208: waveform_sig_loopback =2677;
17209: waveform_sig_loopback =2008;
17210: waveform_sig_loopback =3523;
17211: waveform_sig_loopback =2603;
17212: waveform_sig_loopback =2089;
17213: waveform_sig_loopback =2764;
17214: waveform_sig_loopback =3393;
17215: waveform_sig_loopback =1423;
17216: waveform_sig_loopback =2284;
17217: waveform_sig_loopback =3896;
17218: waveform_sig_loopback =1438;
17219: waveform_sig_loopback =1375;
17220: waveform_sig_loopback =3778;
17221: waveform_sig_loopback =2326;
17222: waveform_sig_loopback =983;
17223: waveform_sig_loopback =2465;
17224: waveform_sig_loopback =3260;
17225: waveform_sig_loopback =957;
17226: waveform_sig_loopback =3589;
17227: waveform_sig_loopback =517;
17228: waveform_sig_loopback =127;
17229: waveform_sig_loopback =4659;
17230: waveform_sig_loopback =1955;
17231: waveform_sig_loopback =802;
17232: waveform_sig_loopback =631;
17233: waveform_sig_loopback =2483;
17234: waveform_sig_loopback =3064;
17235: waveform_sig_loopback =786;
17236: waveform_sig_loopback =844;
17237: waveform_sig_loopback =2241;
17238: waveform_sig_loopback =1125;
17239: waveform_sig_loopback =2160;
17240: waveform_sig_loopback =286;
17241: waveform_sig_loopback =1786;
17242: waveform_sig_loopback =2106;
17243: waveform_sig_loopback =159;
17244: waveform_sig_loopback =1795;
17245: waveform_sig_loopback =936;
17246: waveform_sig_loopback =1301;
17247: waveform_sig_loopback =494;
17248: waveform_sig_loopback =1840;
17249: waveform_sig_loopback =776;
17250: waveform_sig_loopback =188;
17251: waveform_sig_loopback =1672;
17252: waveform_sig_loopback =950;
17253: waveform_sig_loopback =-43;
17254: waveform_sig_loopback =1111;
17255: waveform_sig_loopback =1631;
17256: waveform_sig_loopback =-795;
17257: waveform_sig_loopback =893;
17258: waveform_sig_loopback =1710;
17259: waveform_sig_loopback =-481;
17260: waveform_sig_loopback =-132;
17261: waveform_sig_loopback =1467;
17262: waveform_sig_loopback =728;
17263: waveform_sig_loopback =-1023;
17264: waveform_sig_loopback =471;
17265: waveform_sig_loopback =1700;
17266: waveform_sig_loopback =-1271;
17267: waveform_sig_loopback =1934;
17268: waveform_sig_loopback =-1494;
17269: waveform_sig_loopback =-1827;
17270: waveform_sig_loopback =3100;
17271: waveform_sig_loopback =-181;
17272: waveform_sig_loopback =-1209;
17273: waveform_sig_loopback =-902;
17274: waveform_sig_loopback =440;
17275: waveform_sig_loopback =1148;
17276: waveform_sig_loopback =-1058;
17277: waveform_sig_loopback =-1160;
17278: waveform_sig_loopback =481;
17279: waveform_sig_loopback =-746;
17280: waveform_sig_loopback =95;
17281: waveform_sig_loopback =-1409;
17282: waveform_sig_loopback =-187;
17283: waveform_sig_loopback =-35;
17284: waveform_sig_loopback =-1496;
17285: waveform_sig_loopback =-261;
17286: waveform_sig_loopback =-890;
17287: waveform_sig_loopback =-509;
17288: waveform_sig_loopback =-1643;
17289: waveform_sig_loopback =138;
17290: waveform_sig_loopback =-1211;
17291: waveform_sig_loopback =-1871;
17292: waveform_sig_loopback =132;
17293: waveform_sig_loopback =-1236;
17294: waveform_sig_loopback =-1919;
17295: waveform_sig_loopback =-428;
17296: waveform_sig_loopback =-755;
17297: waveform_sig_loopback =-2386;
17298: waveform_sig_loopback =-940;
17299: waveform_sig_loopback =-412;
17300: waveform_sig_loopback =-2111;
17301: waveform_sig_loopback =-2208;
17302: waveform_sig_loopback =-323;
17303: waveform_sig_loopback =-1094;
17304: waveform_sig_loopback =-3183;
17305: waveform_sig_loopback =-1053;
17306: waveform_sig_loopback =-275;
17307: waveform_sig_loopback =-3316;
17308: waveform_sig_loopback =452;
17309: waveform_sig_loopback =-3793;
17310: waveform_sig_loopback =-3500;
17311: waveform_sig_loopback =1393;
17312: waveform_sig_loopback =-2447;
17313: waveform_sig_loopback =-2906;
17314: waveform_sig_loopback =-2721;
17315: waveform_sig_loopback =-1501;
17316: waveform_sig_loopback =-528;
17317: waveform_sig_loopback =-3191;
17318: waveform_sig_loopback =-2942;
17319: waveform_sig_loopback =-1225;
17320: waveform_sig_loopback =-2768;
17321: waveform_sig_loopback =-1770;
17322: waveform_sig_loopback =-3127;
17323: waveform_sig_loopback =-2100;
17324: waveform_sig_loopback =-1834;
17325: waveform_sig_loopback =-3292;
17326: waveform_sig_loopback =-2290;
17327: waveform_sig_loopback =-2454;
17328: waveform_sig_loopback =-2503;
17329: waveform_sig_loopback =-3559;
17330: waveform_sig_loopback =-1256;
17331: waveform_sig_loopback =-3549;
17332: waveform_sig_loopback =-3367;
17333: waveform_sig_loopback =-1676;
17334: waveform_sig_loopback =-3422;
17335: waveform_sig_loopback =-3285;
17336: waveform_sig_loopback =-2526;
17337: waveform_sig_loopback =-2568;
17338: waveform_sig_loopback =-3997;
17339: waveform_sig_loopback =-2999;
17340: waveform_sig_loopback =-2020;
17341: waveform_sig_loopback =-4034;
17342: waveform_sig_loopback =-4040;
17343: waveform_sig_loopback =-1880;
17344: waveform_sig_loopback =-3120;
17345: waveform_sig_loopback =-4956;
17346: waveform_sig_loopback =-2583;
17347: waveform_sig_loopback =-2329;
17348: waveform_sig_loopback =-5064;
17349: waveform_sig_loopback =-1128;
17350: waveform_sig_loopback =-6006;
17351: waveform_sig_loopback =-4800;
17352: waveform_sig_loopback =-328;
17353: waveform_sig_loopback =-4531;
17354: waveform_sig_loopback =-4333;
17355: waveform_sig_loopback =-4638;
17356: waveform_sig_loopback =-3250;
17357: waveform_sig_loopback =-1981;
17358: waveform_sig_loopback =-5313;
17359: waveform_sig_loopback =-4316;
17360: waveform_sig_loopback =-2985;
17361: waveform_sig_loopback =-4704;
17362: waveform_sig_loopback =-3071;
17363: waveform_sig_loopback =-5151;
17364: waveform_sig_loopback =-3664;
17365: waveform_sig_loopback =-3394;
17366: waveform_sig_loopback =-5216;
17367: waveform_sig_loopback =-3750;
17368: waveform_sig_loopback =-4102;
17369: waveform_sig_loopback =-4450;
17370: waveform_sig_loopback =-4934;
17371: waveform_sig_loopback =-2998;
17372: waveform_sig_loopback =-5303;
17373: waveform_sig_loopback =-4638;
17374: waveform_sig_loopback =-3621;
17375: waveform_sig_loopback =-4982;
17376: waveform_sig_loopback =-4783;
17377: waveform_sig_loopback =-4279;
17378: waveform_sig_loopback =-3940;
17379: waveform_sig_loopback =-5793;
17380: waveform_sig_loopback =-4622;
17381: waveform_sig_loopback =-3313;
17382: waveform_sig_loopback =-5921;
17383: waveform_sig_loopback =-5442;
17384: waveform_sig_loopback =-3289;
17385: waveform_sig_loopback =-5018;
17386: waveform_sig_loopback =-6229;
17387: waveform_sig_loopback =-4017;
17388: waveform_sig_loopback =-4168;
17389: waveform_sig_loopback =-6270;
17390: waveform_sig_loopback =-2783;
17391: waveform_sig_loopback =-7690;
17392: waveform_sig_loopback =-5898;
17393: waveform_sig_loopback =-2211;
17394: waveform_sig_loopback =-5890;
17395: waveform_sig_loopback =-5801;
17396: waveform_sig_loopback =-6337;
17397: waveform_sig_loopback =-4293;
17398: waveform_sig_loopback =-3693;
17399: waveform_sig_loopback =-6953;
17400: waveform_sig_loopback =-5407;
17401: waveform_sig_loopback =-4759;
17402: waveform_sig_loopback =-5926;
17403: waveform_sig_loopback =-4480;
17404: waveform_sig_loopback =-6895;
17405: waveform_sig_loopback =-4673;
17406: waveform_sig_loopback =-4997;
17407: waveform_sig_loopback =-6662;
17408: waveform_sig_loopback =-4940;
17409: waveform_sig_loopback =-5734;
17410: waveform_sig_loopback =-5714;
17411: waveform_sig_loopback =-6076;
17412: waveform_sig_loopback =-4631;
17413: waveform_sig_loopback =-6539;
17414: waveform_sig_loopback =-5960;
17415: waveform_sig_loopback =-5110;
17416: waveform_sig_loopback =-5988;
17417: waveform_sig_loopback =-6411;
17418: waveform_sig_loopback =-5513;
17419: waveform_sig_loopback =-5075;
17420: waveform_sig_loopback =-7400;
17421: waveform_sig_loopback =-5559;
17422: waveform_sig_loopback =-4737;
17423: waveform_sig_loopback =-7362;
17424: waveform_sig_loopback =-6305;
17425: waveform_sig_loopback =-4755;
17426: waveform_sig_loopback =-6206;
17427: waveform_sig_loopback =-7393;
17428: waveform_sig_loopback =-5278;
17429: waveform_sig_loopback =-5381;
17430: waveform_sig_loopback =-7341;
17431: waveform_sig_loopback =-4076;
17432: waveform_sig_loopback =-8989;
17433: waveform_sig_loopback =-6714;
17434: waveform_sig_loopback =-3571;
17435: waveform_sig_loopback =-6901;
17436: waveform_sig_loopback =-7083;
17437: waveform_sig_loopback =-7428;
17438: waveform_sig_loopback =-5090;
17439: waveform_sig_loopback =-5175;
17440: waveform_sig_loopback =-7869;
17441: waveform_sig_loopback =-6399;
17442: waveform_sig_loopback =-6081;
17443: waveform_sig_loopback =-6600;
17444: waveform_sig_loopback =-5840;
17445: waveform_sig_loopback =-7910;
17446: waveform_sig_loopback =-5353;
17447: waveform_sig_loopback =-6465;
17448: waveform_sig_loopback =-7358;
17449: waveform_sig_loopback =-5991;
17450: waveform_sig_loopback =-6842;
17451: waveform_sig_loopback =-6407;
17452: waveform_sig_loopback =-7318;
17453: waveform_sig_loopback =-5488;
17454: waveform_sig_loopback =-7416;
17455: waveform_sig_loopback =-7023;
17456: waveform_sig_loopback =-5839;
17457: waveform_sig_loopback =-7004;
17458: waveform_sig_loopback =-7383;
17459: waveform_sig_loopback =-6095;
17460: waveform_sig_loopback =-6262;
17461: waveform_sig_loopback =-8214;
17462: waveform_sig_loopback =-6129;
17463: waveform_sig_loopback =-5870;
17464: waveform_sig_loopback =-8148;
17465: waveform_sig_loopback =-7050;
17466: waveform_sig_loopback =-5622;
17467: waveform_sig_loopback =-6982;
17468: waveform_sig_loopback =-8279;
17469: waveform_sig_loopback =-5974;
17470: waveform_sig_loopback =-6143;
17471: waveform_sig_loopback =-8072;
17472: waveform_sig_loopback =-4938;
17473: waveform_sig_loopback =-9752;
17474: waveform_sig_loopback =-7329;
17475: waveform_sig_loopback =-4259;
17476: waveform_sig_loopback =-7529;
17477: waveform_sig_loopback =-8057;
17478: waveform_sig_loopback =-7750;
17479: waveform_sig_loopback =-5841;
17480: waveform_sig_loopback =-5980;
17481: waveform_sig_loopback =-8238;
17482: waveform_sig_loopback =-7314;
17483: waveform_sig_loopback =-6501;
17484: waveform_sig_loopback =-7151;
17485: waveform_sig_loopback =-6778;
17486: waveform_sig_loopback =-8046;
17487: waveform_sig_loopback =-6221;
17488: waveform_sig_loopback =-7051;
17489: waveform_sig_loopback =-7622;
17490: waveform_sig_loopback =-6904;
17491: waveform_sig_loopback =-6993;
17492: waveform_sig_loopback =-7150;
17493: waveform_sig_loopback =-7802;
17494: waveform_sig_loopback =-5765;
17495: waveform_sig_loopback =-8261;
17496: waveform_sig_loopback =-7227;
17497: waveform_sig_loopback =-6345;
17498: waveform_sig_loopback =-7513;
17499: waveform_sig_loopback =-7759;
17500: waveform_sig_loopback =-6485;
17501: waveform_sig_loopback =-6743;
17502: waveform_sig_loopback =-8606;
17503: waveform_sig_loopback =-6355;
17504: waveform_sig_loopback =-6474;
17505: waveform_sig_loopback =-8362;
17506: waveform_sig_loopback =-7322;
17507: waveform_sig_loopback =-6152;
17508: waveform_sig_loopback =-7143;
17509: waveform_sig_loopback =-8765;
17510: waveform_sig_loopback =-6117;
17511: waveform_sig_loopback =-6425;
17512: waveform_sig_loopback =-8619;
17513: waveform_sig_loopback =-4846;
17514: waveform_sig_loopback =-10319;
17515: waveform_sig_loopback =-7413;
17516: waveform_sig_loopback =-4250;
17517: waveform_sig_loopback =-8295;
17518: waveform_sig_loopback =-7984;
17519: waveform_sig_loopback =-7802;
17520: waveform_sig_loopback =-6385;
17521: waveform_sig_loopback =-5786;
17522: waveform_sig_loopback =-8821;
17523: waveform_sig_loopback =-7330;
17524: waveform_sig_loopback =-6441;
17525: waveform_sig_loopback =-7744;
17526: waveform_sig_loopback =-6595;
17527: waveform_sig_loopback =-8450;
17528: waveform_sig_loopback =-6252;
17529: waveform_sig_loopback =-6934;
17530: waveform_sig_loopback =-8107;
17531: waveform_sig_loopback =-6906;
17532: waveform_sig_loopback =-7015;
17533: waveform_sig_loopback =-7231;
17534: waveform_sig_loopback =-7747;
17535: waveform_sig_loopback =-6033;
17536: waveform_sig_loopback =-8122;
17537: waveform_sig_loopback =-7188;
17538: waveform_sig_loopback =-6295;
17539: waveform_sig_loopback =-7781;
17540: waveform_sig_loopback =-7553;
17541: waveform_sig_loopback =-6215;
17542: waveform_sig_loopback =-7206;
17543: waveform_sig_loopback =-8130;
17544: waveform_sig_loopback =-6482;
17545: waveform_sig_loopback =-6348;
17546: waveform_sig_loopback =-8142;
17547: waveform_sig_loopback =-7657;
17548: waveform_sig_loopback =-5436;
17549: waveform_sig_loopback =-7374;
17550: waveform_sig_loopback =-8761;
17551: waveform_sig_loopback =-5450;
17552: waveform_sig_loopback =-6855;
17553: waveform_sig_loopback =-7951;
17554: waveform_sig_loopback =-4779;
17555: waveform_sig_loopback =-10591;
17556: waveform_sig_loopback =-6387;
17557: waveform_sig_loopback =-4538;
17558: waveform_sig_loopback =-8060;
17559: waveform_sig_loopback =-7493;
17560: waveform_sig_loopback =-7866;
17561: waveform_sig_loopback =-5750;
17562: waveform_sig_loopback =-5704;
17563: waveform_sig_loopback =-8653;
17564: waveform_sig_loopback =-6633;
17565: waveform_sig_loopback =-6428;
17566: waveform_sig_loopback =-7282;
17567: waveform_sig_loopback =-6114;
17568: waveform_sig_loopback =-8148;
17569: waveform_sig_loopback =-5797;
17570: waveform_sig_loopback =-6686;
17571: waveform_sig_loopback =-7531;
17572: waveform_sig_loopback =-6305;
17573: waveform_sig_loopback =-6708;
17574: waveform_sig_loopback =-7010;
17575: waveform_sig_loopback =-7102;
17576: waveform_sig_loopback =-5370;
17577: waveform_sig_loopback =-8079;
17578: waveform_sig_loopback =-6459;
17579: waveform_sig_loopback =-5899;
17580: waveform_sig_loopback =-7299;
17581: waveform_sig_loopback =-6728;
17582: waveform_sig_loopback =-6214;
17583: waveform_sig_loopback =-6268;
17584: waveform_sig_loopback =-7608;
17585: waveform_sig_loopback =-6146;
17586: waveform_sig_loopback =-5348;
17587: waveform_sig_loopback =-8045;
17588: waveform_sig_loopback =-6634;
17589: waveform_sig_loopback =-4835;
17590: waveform_sig_loopback =-7248;
17591: waveform_sig_loopback =-7486;
17592: waveform_sig_loopback =-5052;
17593: waveform_sig_loopback =-6385;
17594: waveform_sig_loopback =-6869;
17595: waveform_sig_loopback =-4567;
17596: waveform_sig_loopback =-9683;
17597: waveform_sig_loopback =-5603;
17598: waveform_sig_loopback =-4077;
17599: waveform_sig_loopback =-6999;
17600: waveform_sig_loopback =-7071;
17601: waveform_sig_loopback =-7021;
17602: waveform_sig_loopback =-4795;
17603: waveform_sig_loopback =-5087;
17604: waveform_sig_loopback =-7891;
17605: waveform_sig_loopback =-5779;
17606: waveform_sig_loopback =-5715;
17607: waveform_sig_loopback =-6324;
17608: waveform_sig_loopback =-5323;
17609: waveform_sig_loopback =-7482;
17610: waveform_sig_loopback =-4707;
17611: waveform_sig_loopback =-5898;
17612: waveform_sig_loopback =-6820;
17613: waveform_sig_loopback =-5255;
17614: waveform_sig_loopback =-5922;
17615: waveform_sig_loopback =-6138;
17616: waveform_sig_loopback =-5828;
17617: waveform_sig_loopback =-4961;
17618: waveform_sig_loopback =-6787;
17619: waveform_sig_loopback =-5397;
17620: waveform_sig_loopback =-5318;
17621: waveform_sig_loopback =-5814;
17622: waveform_sig_loopback =-6287;
17623: waveform_sig_loopback =-4843;
17624: waveform_sig_loopback =-5236;
17625: waveform_sig_loopback =-7033;
17626: waveform_sig_loopback =-4533;
17627: waveform_sig_loopback =-4764;
17628: waveform_sig_loopback =-6916;
17629: waveform_sig_loopback =-5365;
17630: waveform_sig_loopback =-4033;
17631: waveform_sig_loopback =-5983;
17632: waveform_sig_loopback =-6489;
17633: waveform_sig_loopback =-3939;
17634: waveform_sig_loopback =-5308;
17635: waveform_sig_loopback =-5651;
17636: waveform_sig_loopback =-3584;
17637: waveform_sig_loopback =-8591;
17638: waveform_sig_loopback =-4158;
17639: waveform_sig_loopback =-3125;
17640: waveform_sig_loopback =-5808;
17641: waveform_sig_loopback =-6006;
17642: waveform_sig_loopback =-5792;
17643: waveform_sig_loopback =-3403;
17644: waveform_sig_loopback =-4210;
17645: waveform_sig_loopback =-6539;
17646: waveform_sig_loopback =-4405;
17647: waveform_sig_loopback =-4789;
17648: waveform_sig_loopback =-4749;
17649: waveform_sig_loopback =-4365;
17650: waveform_sig_loopback =-6127;
17651: waveform_sig_loopback =-3179;
17652: waveform_sig_loopback =-5128;
17653: waveform_sig_loopback =-5181;
17654: waveform_sig_loopback =-3988;
17655: waveform_sig_loopback =-4878;
17656: waveform_sig_loopback =-4563;
17657: waveform_sig_loopback =-4713;
17658: waveform_sig_loopback =-3596;
17659: waveform_sig_loopback =-5352;
17660: waveform_sig_loopback =-4365;
17661: waveform_sig_loopback =-3677;
17662: waveform_sig_loopback =-4639;
17663: waveform_sig_loopback =-5009;
17664: waveform_sig_loopback =-3153;
17665: waveform_sig_loopback =-4250;
17666: waveform_sig_loopback =-5461;
17667: waveform_sig_loopback =-3031;
17668: waveform_sig_loopback =-3596;
17669: waveform_sig_loopback =-5389;
17670: waveform_sig_loopback =-3843;
17671: waveform_sig_loopback =-2718;
17672: waveform_sig_loopback =-4559;
17673: waveform_sig_loopback =-4950;
17674: waveform_sig_loopback =-2509;
17675: waveform_sig_loopback =-3833;
17676: waveform_sig_loopback =-4127;
17677: waveform_sig_loopback =-2207;
17678: waveform_sig_loopback =-7003;
17679: waveform_sig_loopback =-2669;
17680: waveform_sig_loopback =-1582;
17681: waveform_sig_loopback =-4260;
17682: waveform_sig_loopback =-4699;
17683: waveform_sig_loopback =-3905;
17684: waveform_sig_loopback =-1979;
17685: waveform_sig_loopback =-2805;
17686: waveform_sig_loopback =-4752;
17687: waveform_sig_loopback =-3061;
17688: waveform_sig_loopback =-3097;
17689: waveform_sig_loopback =-3121;
17690: waveform_sig_loopback =-3079;
17691: waveform_sig_loopback =-4135;
17692: waveform_sig_loopback =-1800;
17693: waveform_sig_loopback =-3645;
17694: waveform_sig_loopback =-3244;
17695: waveform_sig_loopback =-2691;
17696: waveform_sig_loopback =-2984;
17697: waveform_sig_loopback =-3006;
17698: waveform_sig_loopback =-3174;
17699: waveform_sig_loopback =-1686;
17700: waveform_sig_loopback =-4002;
17701: waveform_sig_loopback =-2541;
17702: waveform_sig_loopback =-1877;
17703: waveform_sig_loopback =-3255;
17704: waveform_sig_loopback =-3132;
17705: waveform_sig_loopback =-1478;
17706: waveform_sig_loopback =-2669;
17707: waveform_sig_loopback =-3586;
17708: waveform_sig_loopback =-1413;
17709: waveform_sig_loopback =-2010;
17710: waveform_sig_loopback =-3568;
17711: waveform_sig_loopback =-2082;
17712: waveform_sig_loopback =-1136;
17713: waveform_sig_loopback =-2776;
17714: waveform_sig_loopback =-3280;
17715: waveform_sig_loopback =-622;
17716: waveform_sig_loopback =-2173;
17717: waveform_sig_loopback =-2533;
17718: waveform_sig_loopback =-329;
17719: waveform_sig_loopback =-5383;
17720: waveform_sig_loopback =-805;
17721: waveform_sig_loopback =276;
17722: waveform_sig_loopback =-2855;
17723: waveform_sig_loopback =-2758;
17724: waveform_sig_loopback =-2063;
17725: waveform_sig_loopback =-403;
17726: waveform_sig_loopback =-869;
17727: waveform_sig_loopback =-3187;
17728: waveform_sig_loopback =-1225;
17729: waveform_sig_loopback =-1148;
17730: waveform_sig_loopback =-1443;
17731: waveform_sig_loopback =-1355;
17732: waveform_sig_loopback =-2190;
17733: waveform_sig_loopback =-136;
17734: waveform_sig_loopback =-1746;
17735: waveform_sig_loopback =-1414;
17736: waveform_sig_loopback =-1000;
17737: waveform_sig_loopback =-974;
17738: waveform_sig_loopback =-1353;
17739: waveform_sig_loopback =-1275;
17740: waveform_sig_loopback =188;
17741: waveform_sig_loopback =-2298;
17742: waveform_sig_loopback =-529;
17743: waveform_sig_loopback =-59;
17744: waveform_sig_loopback =-1634;
17745: waveform_sig_loopback =-940;
17746: waveform_sig_loopback =290;
17747: waveform_sig_loopback =-1167;
17748: waveform_sig_loopback =-1378;
17749: waveform_sig_loopback =413;
17750: waveform_sig_loopback =-173;
17751: waveform_sig_loopback =-1814;
17752: waveform_sig_loopback =-200;
17753: waveform_sig_loopback =1000;
17754: waveform_sig_loopback =-1171;
17755: waveform_sig_loopback =-1494;
17756: waveform_sig_loopback =1549;
17757: waveform_sig_loopback =-522;
17758: waveform_sig_loopback =-550;
17759: waveform_sig_loopback =1513;
17760: waveform_sig_loopback =-3736;
17761: waveform_sig_loopback =1429;
17762: waveform_sig_loopback =2006;
17763: waveform_sig_loopback =-1212;
17764: waveform_sig_loopback =-566;
17765: waveform_sig_loopback =-296;
17766: waveform_sig_loopback =1452;
17767: waveform_sig_loopback =1205;
17768: waveform_sig_loopback =-1636;
17769: waveform_sig_loopback =967;
17770: waveform_sig_loopback =632;
17771: waveform_sig_loopback =242;
17772: waveform_sig_loopback =845;
17773: waveform_sig_loopback =-488;
17774: waveform_sig_loopback =1789;
17775: waveform_sig_loopback =228;
17776: waveform_sig_loopback =342;
17777: waveform_sig_loopback =997;
17778: waveform_sig_loopback =944;
17779: waveform_sig_loopback =240;
17780: waveform_sig_loopback =1017;
17781: waveform_sig_loopback =1853;
17782: waveform_sig_loopback =-608;
17783: waveform_sig_loopback =1755;
17784: waveform_sig_loopback =1453;
17785: waveform_sig_loopback =373;
17786: waveform_sig_loopback =1028;
17787: waveform_sig_loopback =2022;
17788: waveform_sig_loopback =901;
17789: waveform_sig_loopback =373;
17790: waveform_sig_loopback =2324;
17791: waveform_sig_loopback =1772;
17792: waveform_sig_loopback =15;
17793: waveform_sig_loopback =1677;
17794: waveform_sig_loopback =2997;
17795: waveform_sig_loopback =475;
17796: waveform_sig_loopback =507;
17797: waveform_sig_loopback =3654;
17798: waveform_sig_loopback =820;
17799: waveform_sig_loopback =1884;
17800: waveform_sig_loopback =3088;
17801: waveform_sig_loopback =-2032;
17802: waveform_sig_loopback =3977;
17803: waveform_sig_loopback =3248;
17804: waveform_sig_loopback =927;
17805: waveform_sig_loopback =1358;
17806: waveform_sig_loopback =1254;
17807: waveform_sig_loopback =3828;
17808: waveform_sig_loopback =2640;
17809: waveform_sig_loopback =246;
17810: waveform_sig_loopback =3196;
17811: waveform_sig_loopback =2068;
17812: waveform_sig_loopback =2417;
17813: waveform_sig_loopback =2532;
17814: waveform_sig_loopback =1252;
17815: waveform_sig_loopback =3931;
17816: waveform_sig_loopback =1829;
17817: waveform_sig_loopback =2193;
17818: waveform_sig_loopback =2979;
17819: waveform_sig_loopback =2662;
17820: waveform_sig_loopback =2114;
17821: waveform_sig_loopback =3015;
17822: waveform_sig_loopback =3395;
17823: waveform_sig_loopback =1351;
17824: waveform_sig_loopback =3766;
17825: waveform_sig_loopback =3013;
17826: waveform_sig_loopback =2406;
17827: waveform_sig_loopback =2696;
17828: waveform_sig_loopback =3840;
17829: waveform_sig_loopback =2884;
17830: waveform_sig_loopback =1878;
17831: waveform_sig_loopback =4352;
17832: waveform_sig_loopback =3492;
17833: waveform_sig_loopback =1637;
17834: waveform_sig_loopback =3784;
17835: waveform_sig_loopback =4606;
17836: waveform_sig_loopback =2101;
17837: waveform_sig_loopback =2634;
17838: waveform_sig_loopback =5228;
17839: waveform_sig_loopback =2488;
17840: waveform_sig_loopback =4052;
17841: waveform_sig_loopback =4300;
17842: waveform_sig_loopback =45;
17843: waveform_sig_loopback =5849;
17844: waveform_sig_loopback =4647;
17845: waveform_sig_loopback =3092;
17846: waveform_sig_loopback =2701;
17847: waveform_sig_loopback =3260;
17848: waveform_sig_loopback =5765;
17849: waveform_sig_loopback =3879;
17850: waveform_sig_loopback =2325;
17851: waveform_sig_loopback =4796;
17852: waveform_sig_loopback =3658;
17853: waveform_sig_loopback =4461;
17854: waveform_sig_loopback =3900;
17855: waveform_sig_loopback =3111;
17856: waveform_sig_loopback =5693;
17857: waveform_sig_loopback =3282;
17858: waveform_sig_loopback =4080;
17859: waveform_sig_loopback =4565;
17860: waveform_sig_loopback =4244;
17861: waveform_sig_loopback =3815;
17862: waveform_sig_loopback =4764;
17863: waveform_sig_loopback =4851;
17864: waveform_sig_loopback =3214;
17865: waveform_sig_loopback =5254;
17866: waveform_sig_loopback =4535;
17867: waveform_sig_loopback =4272;
17868: waveform_sig_loopback =3989;
17869: waveform_sig_loopback =5732;
17870: waveform_sig_loopback =4347;
17871: waveform_sig_loopback =3216;
17872: waveform_sig_loopback =6436;
17873: waveform_sig_loopback =4581;
17874: waveform_sig_loopback =3306;
17875: waveform_sig_loopback =5501;
17876: waveform_sig_loopback =5699;
17877: waveform_sig_loopback =4120;
17878: waveform_sig_loopback =4021;
17879: waveform_sig_loopback =6533;
17880: waveform_sig_loopback =4120;
17881: waveform_sig_loopback =5582;
17882: waveform_sig_loopback =5800;
17883: waveform_sig_loopback =1464;
17884: waveform_sig_loopback =7264;
17885: waveform_sig_loopback =6375;
17886: waveform_sig_loopback =4380;
17887: waveform_sig_loopback =4021;
17888: waveform_sig_loopback =4978;
17889: waveform_sig_loopback =7097;
17890: waveform_sig_loopback =5265;
17891: waveform_sig_loopback =3829;
17892: waveform_sig_loopback =6150;
17893: waveform_sig_loopback =5136;
17894: waveform_sig_loopback =5931;
17895: waveform_sig_loopback =4992;
17896: waveform_sig_loopback =4770;
17897: waveform_sig_loopback =7076;
17898: waveform_sig_loopback =4377;
17899: waveform_sig_loopback =5724;
17900: waveform_sig_loopback =5776;
17901: waveform_sig_loopback =5601;
17902: waveform_sig_loopback =5325;
17903: waveform_sig_loopback =5737;
17904: waveform_sig_loopback =6402;
17905: waveform_sig_loopback =4556;
17906: waveform_sig_loopback =6302;
17907: waveform_sig_loopback =6194;
17908: waveform_sig_loopback =5198;
17909: waveform_sig_loopback =5512;
17910: waveform_sig_loopback =7070;
17911: waveform_sig_loopback =5108;
17912: waveform_sig_loopback =5032;
17913: waveform_sig_loopback =7471;
17914: waveform_sig_loopback =5643;
17915: waveform_sig_loopback =4755;
17916: waveform_sig_loopback =6730;
17917: waveform_sig_loopback =6926;
17918: waveform_sig_loopback =5119;
17919: waveform_sig_loopback =5218;
17920: waveform_sig_loopback =7935;
17921: waveform_sig_loopback =5294;
17922: waveform_sig_loopback =6545;
17923: waveform_sig_loopback =6893;
17924: waveform_sig_loopback =2835;
17925: waveform_sig_loopback =8493;
17926: waveform_sig_loopback =7386;
17927: waveform_sig_loopback =5284;
17928: waveform_sig_loopback =5284;
17929: waveform_sig_loopback =6322;
17930: waveform_sig_loopback =7828;
17931: waveform_sig_loopback =6439;
17932: waveform_sig_loopback =5044;
17933: waveform_sig_loopback =7025;
17934: waveform_sig_loopback =6417;
17935: waveform_sig_loopback =6753;
17936: waveform_sig_loopback =6095;
17937: waveform_sig_loopback =6130;
17938: waveform_sig_loopback =7611;
17939: waveform_sig_loopback =5673;
17940: waveform_sig_loopback =6754;
17941: waveform_sig_loopback =6503;
17942: waveform_sig_loopback =6886;
17943: waveform_sig_loopback =5978;
17944: waveform_sig_loopback =6951;
17945: waveform_sig_loopback =7384;
17946: waveform_sig_loopback =5162;
17947: waveform_sig_loopback =7549;
17948: waveform_sig_loopback =7046;
17949: waveform_sig_loopback =5908;
17950: waveform_sig_loopback =6701;
17951: waveform_sig_loopback =7804;
17952: waveform_sig_loopback =5974;
17953: waveform_sig_loopback =6121;
17954: waveform_sig_loopback =8153;
17955: waveform_sig_loopback =6527;
17956: waveform_sig_loopback =5666;
17957: waveform_sig_loopback =7506;
17958: waveform_sig_loopback =7806;
17959: waveform_sig_loopback =5869;
17960: waveform_sig_loopback =6014;
17961: waveform_sig_loopback =8940;
17962: waveform_sig_loopback =5797;
17963: waveform_sig_loopback =7469;
17964: waveform_sig_loopback =7625;
17965: waveform_sig_loopback =3352;
17966: waveform_sig_loopback =9574;
17967: waveform_sig_loopback =8008;
17968: waveform_sig_loopback =5704;
17969: waveform_sig_loopback =6339;
17970: waveform_sig_loopback =6838;
17971: waveform_sig_loopback =8496;
17972: waveform_sig_loopback =7310;
17973: waveform_sig_loopback =5316;
17974: waveform_sig_loopback =7990;
17975: waveform_sig_loopback =6975;
17976: waveform_sig_loopback =7171;
17977: waveform_sig_loopback =7002;
17978: waveform_sig_loopback =6451;
17979: waveform_sig_loopback =8292;
17980: waveform_sig_loopback =6406;
17981: waveform_sig_loopback =7023;
17982: waveform_sig_loopback =7354;
17983: waveform_sig_loopback =7297;
17984: waveform_sig_loopback =6419;
17985: waveform_sig_loopback =7720;
17986: waveform_sig_loopback =7598;
17987: waveform_sig_loopback =5832;
17988: waveform_sig_loopback =8097;
17989: waveform_sig_loopback =7422;
17990: waveform_sig_loopback =6309;
17991: waveform_sig_loopback =7341;
17992: waveform_sig_loopback =8131;
17993: waveform_sig_loopback =6251;
17994: waveform_sig_loopback =6834;
17995: waveform_sig_loopback =8250;
17996: waveform_sig_loopback =7101;
17997: waveform_sig_loopback =5979;
17998: waveform_sig_loopback =7759;
17999: waveform_sig_loopback =8559;
18000: waveform_sig_loopback =5712;
18001: waveform_sig_loopback =6646;
18002: waveform_sig_loopback =9404;
18003: waveform_sig_loopback =5614;
18004: waveform_sig_loopback =8471;
18005: waveform_sig_loopback =7277;
18006: waveform_sig_loopback =3755;
18007: waveform_sig_loopback =10309;
18008: waveform_sig_loopback =7593;
18009: waveform_sig_loopback =6374;
18010: waveform_sig_loopback =6400;
18011: waveform_sig_loopback =6918;
18012: waveform_sig_loopback =9146;
18013: waveform_sig_loopback =6986;
18014: waveform_sig_loopback =5705;
18015: waveform_sig_loopback =8275;
18016: waveform_sig_loopback =6830;
18017: waveform_sig_loopback =7596;
18018: waveform_sig_loopback =6917;
18019: waveform_sig_loopback =6604;
18020: waveform_sig_loopback =8498;
18021: waveform_sig_loopback =6331;
18022: waveform_sig_loopback =7198;
18023: waveform_sig_loopback =7419;
18024: waveform_sig_loopback =7348;
18025: waveform_sig_loopback =6337;
18026: waveform_sig_loopback =8028;
18027: waveform_sig_loopback =7349;
18028: waveform_sig_loopback =5861;
18029: waveform_sig_loopback =8390;
18030: waveform_sig_loopback =6953;
18031: waveform_sig_loopback =6652;
18032: waveform_sig_loopback =7217;
18033: waveform_sig_loopback =7887;
18034: waveform_sig_loopback =6586;
18035: waveform_sig_loopback =6408;
18036: waveform_sig_loopback =8452;
18037: waveform_sig_loopback =7029;
18038: waveform_sig_loopback =5524;
18039: waveform_sig_loopback =8221;
18040: waveform_sig_loopback =8007;
18041: waveform_sig_loopback =5468;
18042: waveform_sig_loopback =6997;
18043: waveform_sig_loopback =8671;
18044: waveform_sig_loopback =5706;
18045: waveform_sig_loopback =8344;
18046: waveform_sig_loopback =6586;
18047: waveform_sig_loopback =4092;
18048: waveform_sig_loopback =9833;
18049: waveform_sig_loopback =7296;
18050: waveform_sig_loopback =6266;
18051: waveform_sig_loopback =5896;
18052: waveform_sig_loopback =6885;
18053: waveform_sig_loopback =8846;
18054: waveform_sig_loopback =6453;
18055: waveform_sig_loopback =5521;
18056: waveform_sig_loopback =7988;
18057: waveform_sig_loopback =6308;
18058: waveform_sig_loopback =7532;
18059: waveform_sig_loopback =6308;
18060: waveform_sig_loopback =6296;
18061: waveform_sig_loopback =8253;
18062: waveform_sig_loopback =5699;
18063: waveform_sig_loopback =6934;
18064: waveform_sig_loopback =7058;
18065: waveform_sig_loopback =6658;
18066: waveform_sig_loopback =6172;
18067: waveform_sig_loopback =7607;
18068: waveform_sig_loopback =6558;
18069: waveform_sig_loopback =5850;
18070: waveform_sig_loopback =7551;
18071: waveform_sig_loopback =6577;
18072: waveform_sig_loopback =6278;
18073: waveform_sig_loopback =6354;
18074: waveform_sig_loopback =7783;
18075: waveform_sig_loopback =5715;
18076: waveform_sig_loopback =5811;
18077: waveform_sig_loopback =8190;
18078: waveform_sig_loopback =5960;
18079: waveform_sig_loopback =5189;
18080: waveform_sig_loopback =7670;
18081: waveform_sig_loopback =7079;
18082: waveform_sig_loopback =5105;
18083: waveform_sig_loopback =6238;
18084: waveform_sig_loopback =7928;
18085: waveform_sig_loopback =5146;
18086: waveform_sig_loopback =7606;
18087: waveform_sig_loopback =5778;
18088: waveform_sig_loopback =3537;
18089: waveform_sig_loopback =9097;
18090: waveform_sig_loopback =6576;
18091: waveform_sig_loopback =5413;
18092: waveform_sig_loopback =5104;
18093: waveform_sig_loopback =6303;
18094: waveform_sig_loopback =8008;
18095: waveform_sig_loopback =5513;
18096: waveform_sig_loopback =4966;
18097: waveform_sig_loopback =7125;
18098: waveform_sig_loopback =5418;
18099: waveform_sig_loopback =6914;
18100: waveform_sig_loopback =5193;
18101: waveform_sig_loopback =5754;
18102: waveform_sig_loopback =7336;
18103: waveform_sig_loopback =4522;
18104: waveform_sig_loopback =6509;
18105: waveform_sig_loopback =5860;
18106: waveform_sig_loopback =5761;
18107: waveform_sig_loopback =5509;
18108: waveform_sig_loopback =6256;
18109: waveform_sig_loopback =5964;
18110: waveform_sig_loopback =4758;
18111: waveform_sig_loopback =6408;
18112: waveform_sig_loopback =5991;
18113: waveform_sig_loopback =4827;
18114: waveform_sig_loopback =5769;
18115: waveform_sig_loopback =6667;
18116: waveform_sig_loopback =4415;
18117: waveform_sig_loopback =5252;
18118: waveform_sig_loopback =6926;
18119: waveform_sig_loopback =4878;
18120: waveform_sig_loopback =4260;
18121: waveform_sig_loopback =6641;
18122: waveform_sig_loopback =5930;
18123: waveform_sig_loopback =4033;
18124: waveform_sig_loopback =5263;
18125: waveform_sig_loopback =6769;
18126: waveform_sig_loopback =4119;
18127: waveform_sig_loopback =6446;
18128: waveform_sig_loopback =4538;
18129: waveform_sig_loopback =2640;
18130: waveform_sig_loopback =7817;
18131: waveform_sig_loopback =5584;
18132: waveform_sig_loopback =4076;
18133: waveform_sig_loopback =3956;
18134: waveform_sig_loopback =5447;
18135: waveform_sig_loopback =6471;
18136: waveform_sig_loopback =4486;
18137: waveform_sig_loopback =3814;
18138: waveform_sig_loopback =5664;
18139: waveform_sig_loopback =4533;
18140: waveform_sig_loopback =5414;
18141: waveform_sig_loopback =3894;
18142: waveform_sig_loopback =4822;
18143: waveform_sig_loopback =5681;
18144: waveform_sig_loopback =3527;
18145: waveform_sig_loopback =5157;
18146: waveform_sig_loopback =4325;
18147: waveform_sig_loopback =4812;
18148: waveform_sig_loopback =3894;
18149: waveform_sig_loopback =5151;
18150: waveform_sig_loopback =4625;
18151: waveform_sig_loopback =3196;
18152: waveform_sig_loopback =5359;
18153: waveform_sig_loopback =4460;
18154: waveform_sig_loopback =3335;
18155: waveform_sig_loopback =4622;
18156: waveform_sig_loopback =5150;
18157: waveform_sig_loopback =2953;
18158: waveform_sig_loopback =4067;
18159: waveform_sig_loopback =5349;
18160: waveform_sig_loopback =3448;
18161: waveform_sig_loopback =3021;
18162: waveform_sig_loopback =5011;
18163: waveform_sig_loopback =4641;
18164: waveform_sig_loopback =2476;
18165: waveform_sig_loopback =3735;
18166: waveform_sig_loopback =5548;
18167: waveform_sig_loopback =2393;
18168: waveform_sig_loopback =5154;
18169: waveform_sig_loopback =2964;
18170: waveform_sig_loopback =1024;
18171: waveform_sig_loopback =6584;
18172: waveform_sig_loopback =3916;
18173: waveform_sig_loopback =2410;
18174: waveform_sig_loopback =2674;
18175: waveform_sig_loopback =3803;
18176: waveform_sig_loopback =4894;
18177: waveform_sig_loopback =3107;
18178: waveform_sig_loopback =2020;
18179: waveform_sig_loopback =4309;
18180: waveform_sig_loopback =2997;
18181: waveform_sig_loopback =3629;
18182: waveform_sig_loopback =2640;
18183: waveform_sig_loopback =3123;
18184: waveform_sig_loopback =4004;
18185: waveform_sig_loopback =2213;
18186: waveform_sig_loopback =3311;
18187: waveform_sig_loopback =2949;
18188: waveform_sig_loopback =3199;
18189: waveform_sig_loopback =2068;
18190: waveform_sig_loopback =3904;
18191: waveform_sig_loopback =2678;
18192: waveform_sig_loopback =1656;
18193: waveform_sig_loopback =3958;
18194: waveform_sig_loopback =2532;
18195: waveform_sig_loopback =1846;
18196: waveform_sig_loopback =3071;
18197: waveform_sig_loopback =3291;
18198: waveform_sig_loopback =1450;
18199: waveform_sig_loopback =2423;
18200: waveform_sig_loopback =3570;
18201: waveform_sig_loopback =1855;
18202: waveform_sig_loopback =1294;
18203: waveform_sig_loopback =3384;
18204: waveform_sig_loopback =2964;
18205: waveform_sig_loopback =583;
18206: waveform_sig_loopback =2336;
18207: waveform_sig_loopback =3823;
18208: waveform_sig_loopback =358;
18209: waveform_sig_loopback =3871;
18210: waveform_sig_loopback =816;
18211: waveform_sig_loopback =-525;
18212: waveform_sig_loopback =5206;
18213: waveform_sig_loopback =1709;
18214: waveform_sig_loopback =842;
18215: waveform_sig_loopback =1036;
18216: waveform_sig_loopback =1813;
18217: waveform_sig_loopback =3488;
18218: waveform_sig_loopback =970;
18219: waveform_sig_loopback =302;
18220: waveform_sig_loopback =2752;
18221: waveform_sig_loopback =904;
18222: waveform_sig_loopback =2012;
18223: waveform_sig_loopback =830;
18224: waveform_sig_loopback =982;
18225: waveform_sig_loopback =2472;
18226: waveform_sig_loopback =409;
18227: waveform_sig_loopback =1350;
18228: waveform_sig_loopback =1264;
18229: waveform_sig_loopback =1072;
18230: waveform_sig_loopback =549;
18231: waveform_sig_loopback =2163;
18232: waveform_sig_loopback =413;
18233: waveform_sig_loopback =123;
18234: waveform_sig_loopback =2196;
18235: waveform_sig_loopback =507;
18236: waveform_sig_loopback =138;
18237: waveform_sig_loopback =1134;
18238: waveform_sig_loopback =1415;
18239: waveform_sig_loopback =-299;
18240: waveform_sig_loopback =370;
18241: waveform_sig_loopback =1834;
18242: waveform_sig_loopback =4;
18243: waveform_sig_loopback =-729;
18244: waveform_sig_loopback =1684;
18245: waveform_sig_loopback =943;
18246: waveform_sig_loopback =-1352;
18247: waveform_sig_loopback =751;
18248: waveform_sig_loopback =1630;
18249: waveform_sig_loopback =-1454;
18250: waveform_sig_loopback =2368;
18251: waveform_sig_loopback =-1711;
18252: waveform_sig_loopback =-1975;
18253: waveform_sig_loopback =3354;
18254: waveform_sig_loopback =-613;
18255: waveform_sig_loopback =-662;
18256: waveform_sig_loopback =-1145;
18257: waveform_sig_loopback =110;
18258: waveform_sig_loopback =1839;
18259: waveform_sig_loopback =-1590;
18260: waveform_sig_loopback =-1101;
18261: waveform_sig_loopback =789;
18262: waveform_sig_loopback =-1221;
18263: waveform_sig_loopback =553;
18264: waveform_sig_loopback =-1634;
18265: waveform_sig_loopback =-359;
18266: waveform_sig_loopback =520;
18267: waveform_sig_loopback =-1967;
18268: waveform_sig_loopback =-116;
18269: waveform_sig_loopback =-737;
18270: waveform_sig_loopback =-798;
18271: waveform_sig_loopback =-1449;
18272: waveform_sig_loopback =184;
18273: waveform_sig_loopback =-1412;
18274: waveform_sig_loopback =-1595;
18275: waveform_sig_loopback =57;
18276: waveform_sig_loopback =-1493;
18277: waveform_sig_loopback =-1509;
18278: waveform_sig_loopback =-861;
18279: waveform_sig_loopback =-506;
18280: waveform_sig_loopback =-2152;
18281: waveform_sig_loopback =-1567;
18282: waveform_sig_loopback =200;
18283: waveform_sig_loopback =-2280;
18284: waveform_sig_loopback =-2531;
18285: waveform_sig_loopback =251;
18286: waveform_sig_loopback =-1494;
18287: waveform_sig_loopback =-3057;
18288: waveform_sig_loopback =-943;
18289: waveform_sig_loopback =-651;
18290: waveform_sig_loopback =-2921;
18291: waveform_sig_loopback =145;
18292: waveform_sig_loopback =-3761;
18293: waveform_sig_loopback =-3227;
18294: waveform_sig_loopback =952;
18295: waveform_sig_loopback =-2183;
18296: waveform_sig_loopback =-2620;
18297: waveform_sig_loopback =-3298;
18298: waveform_sig_loopback =-1239;
18299: waveform_sig_loopback =-462;
18300: waveform_sig_loopback =-3359;
18301: waveform_sig_loopback =-2672;
18302: waveform_sig_loopback =-1480;
18303: waveform_sig_loopback =-2751;
18304: waveform_sig_loopback =-1415;
18305: waveform_sig_loopback =-3612;
18306: waveform_sig_loopback =-1891;
18307: waveform_sig_loopback =-1649;
18308: waveform_sig_loopback =-3670;
18309: waveform_sig_loopback =-1933;
18310: waveform_sig_loopback =-2680;
18311: waveform_sig_loopback =-2629;
18312: waveform_sig_loopback =-3192;
18313: waveform_sig_loopback =-1664;
18314: waveform_sig_loopback =-3410;
18315: waveform_sig_loopback =-3169;
18316: waveform_sig_loopback =-2087;
18317: waveform_sig_loopback =-3059;
18318: waveform_sig_loopback =-3395;
18319: waveform_sig_loopback =-2852;
18320: waveform_sig_loopback =-1897;
18321: waveform_sig_loopback =-4500;
18322: waveform_sig_loopback =-3016;
18323: waveform_sig_loopback =-1564;
18324: waveform_sig_loopback =-4539;
18325: waveform_sig_loopback =-3746;
18326: waveform_sig_loopback =-1935;
18327: waveform_sig_loopback =-3280;
18328: waveform_sig_loopback =-4535;
18329: waveform_sig_loopback =-3059;
18330: waveform_sig_loopback =-2133;
18331: waveform_sig_loopback =-4791;
18332: waveform_sig_loopback =-1679;
18333: waveform_sig_loopback =-5420;
18334: waveform_sig_loopback =-5073;
18335: waveform_sig_loopback =-702;
18336: waveform_sig_loopback =-3933;
18337: waveform_sig_loopback =-4589;
18338: waveform_sig_loopback =-4753;
18339: waveform_sig_loopback =-2963;
18340: waveform_sig_loopback =-2361;
18341: waveform_sig_loopback =-4968;
18342: waveform_sig_loopback =-4399;
18343: waveform_sig_loopback =-3220;
18344: waveform_sig_loopback =-4320;
18345: waveform_sig_loopback =-3283;
18346: waveform_sig_loopback =-5228;
18347: waveform_sig_loopback =-3442;
18348: waveform_sig_loopback =-3538;
18349: waveform_sig_loopback =-5237;
18350: waveform_sig_loopback =-3522;
18351: waveform_sig_loopback =-4463;
18352: waveform_sig_loopback =-4221;
18353: waveform_sig_loopback =-4773;
18354: waveform_sig_loopback =-3497;
18355: waveform_sig_loopback =-4798;
18356: waveform_sig_loopback =-4996;
18357: waveform_sig_loopback =-3647;
18358: waveform_sig_loopback =-4430;
18359: waveform_sig_loopback =-5502;
18360: waveform_sig_loopback =-3899;
18361: waveform_sig_loopback =-3817;
18362: waveform_sig_loopback =-6247;
18363: waveform_sig_loopback =-4051;
18364: waveform_sig_loopback =-3696;
18365: waveform_sig_loopback =-5801;
18366: waveform_sig_loopback =-5248;
18367: waveform_sig_loopback =-3739;
18368: waveform_sig_loopback =-4489;
18369: waveform_sig_loopback =-6481;
18370: waveform_sig_loopback =-4321;
18371: waveform_sig_loopback =-3636;
18372: waveform_sig_loopback =-6613;
18373: waveform_sig_loopback =-2850;
18374: waveform_sig_loopback =-7304;
18375: waveform_sig_loopback =-6323;
18376: waveform_sig_loopback =-2117;
18377: waveform_sig_loopback =-5678;
18378: waveform_sig_loopback =-6006;
18379: waveform_sig_loopback =-6147;
18380: waveform_sig_loopback =-4336;
18381: waveform_sig_loopback =-4007;
18382: waveform_sig_loopback =-6390;
18383: waveform_sig_loopback =-5800;
18384: waveform_sig_loopback =-4724;
18385: waveform_sig_loopback =-5536;
18386: waveform_sig_loopback =-5067;
18387: waveform_sig_loopback =-6372;
18388: waveform_sig_loopback =-4771;
18389: waveform_sig_loopback =-5247;
18390: waveform_sig_loopback =-6178;
18391: waveform_sig_loopback =-5261;
18392: waveform_sig_loopback =-5621;
18393: waveform_sig_loopback =-5415;
18394: waveform_sig_loopback =-6598;
18395: waveform_sig_loopback =-4321;
18396: waveform_sig_loopback =-6491;
18397: waveform_sig_loopback =-6380;
18398: waveform_sig_loopback =-4634;
18399: waveform_sig_loopback =-6277;
18400: waveform_sig_loopback =-6466;
18401: waveform_sig_loopback =-5225;
18402: waveform_sig_loopback =-5444;
18403: waveform_sig_loopback =-7158;
18404: waveform_sig_loopback =-5513;
18405: waveform_sig_loopback =-4965;
18406: waveform_sig_loopback =-7050;
18407: waveform_sig_loopback =-6566;
18408: waveform_sig_loopback =-4791;
18409: waveform_sig_loopback =-5871;
18410: waveform_sig_loopback =-7749;
18411: waveform_sig_loopback =-5367;
18412: waveform_sig_loopback =-4951;
18413: waveform_sig_loopback =-7863;
18414: waveform_sig_loopback =-3968;
18415: waveform_sig_loopback =-8632;
18416: waveform_sig_loopback =-7405;
18417: waveform_sig_loopback =-3132;
18418: waveform_sig_loopback =-7078;
18419: waveform_sig_loopback =-7123;
18420: waveform_sig_loopback =-7042;
18421: waveform_sig_loopback =-5768;
18422: waveform_sig_loopback =-4798;
18423: waveform_sig_loopback =-7646;
18424: waveform_sig_loopback =-7019;
18425: waveform_sig_loopback =-5472;
18426: waveform_sig_loopback =-6949;
18427: waveform_sig_loopback =-5907;
18428: waveform_sig_loopback =-7367;
18429: waveform_sig_loopback =-6054;
18430: waveform_sig_loopback =-6003;
18431: waveform_sig_loopback =-7382;
18432: waveform_sig_loopback =-6320;
18433: waveform_sig_loopback =-6388;
18434: waveform_sig_loopback =-6725;
18435: waveform_sig_loopback =-7284;
18436: waveform_sig_loopback =-5247;
18437: waveform_sig_loopback =-7720;
18438: waveform_sig_loopback =-6921;
18439: waveform_sig_loopback =-5723;
18440: waveform_sig_loopback =-7248;
18441: waveform_sig_loopback =-7187;
18442: waveform_sig_loopback =-6176;
18443: waveform_sig_loopback =-6357;
18444: waveform_sig_loopback =-7934;
18445: waveform_sig_loopback =-6403;
18446: waveform_sig_loopback =-5795;
18447: waveform_sig_loopback =-7851;
18448: waveform_sig_loopback =-7501;
18449: waveform_sig_loopback =-5384;
18450: waveform_sig_loopback =-6796;
18451: waveform_sig_loopback =-8694;
18452: waveform_sig_loopback =-5738;
18453: waveform_sig_loopback =-6089;
18454: waveform_sig_loopback =-8408;
18455: waveform_sig_loopback =-4542;
18456: waveform_sig_loopback =-9918;
18457: waveform_sig_loopback =-7420;
18458: waveform_sig_loopback =-4015;
18459: waveform_sig_loopback =-8058;
18460: waveform_sig_loopback =-7476;
18461: waveform_sig_loopback =-7950;
18462: waveform_sig_loopback =-6247;
18463: waveform_sig_loopback =-5406;
18464: waveform_sig_loopback =-8723;
18465: waveform_sig_loopback =-7128;
18466: waveform_sig_loopback =-6326;
18467: waveform_sig_loopback =-7749;
18468: waveform_sig_loopback =-6139;
18469: waveform_sig_loopback =-8341;
18470: waveform_sig_loopback =-6403;
18471: waveform_sig_loopback =-6596;
18472: waveform_sig_loopback =-8118;
18473: waveform_sig_loopback =-6540;
18474: waveform_sig_loopback =-7132;
18475: waveform_sig_loopback =-7323;
18476: waveform_sig_loopback =-7559;
18477: waveform_sig_loopback =-5904;
18478: waveform_sig_loopback =-8294;
18479: waveform_sig_loopback =-7238;
18480: waveform_sig_loopback =-6292;
18481: waveform_sig_loopback =-7710;
18482: waveform_sig_loopback =-7499;
18483: waveform_sig_loopback =-6749;
18484: waveform_sig_loopback =-6699;
18485: waveform_sig_loopback =-8334;
18486: waveform_sig_loopback =-6960;
18487: waveform_sig_loopback =-5936;
18488: waveform_sig_loopback =-8496;
18489: waveform_sig_loopback =-7816;
18490: waveform_sig_loopback =-5492;
18491: waveform_sig_loopback =-7611;
18492: waveform_sig_loopback =-8634;
18493: waveform_sig_loopback =-6017;
18494: waveform_sig_loopback =-6820;
18495: waveform_sig_loopback =-8145;
18496: waveform_sig_loopback =-5168;
18497: waveform_sig_loopback =-10249;
18498: waveform_sig_loopback =-7281;
18499: waveform_sig_loopback =-4758;
18500: waveform_sig_loopback =-7855;
18501: waveform_sig_loopback =-7898;
18502: waveform_sig_loopback =-8390;
18503: waveform_sig_loopback =-5984;
18504: waveform_sig_loopback =-5843;
18505: waveform_sig_loopback =-8905;
18506: waveform_sig_loopback =-7193;
18507: waveform_sig_loopback =-6715;
18508: waveform_sig_loopback =-7586;
18509: waveform_sig_loopback =-6406;
18510: waveform_sig_loopback =-8697;
18511: waveform_sig_loopback =-6143;
18512: waveform_sig_loopback =-6919;
18513: waveform_sig_loopback =-8243;
18514: waveform_sig_loopback =-6535;
18515: waveform_sig_loopback =-7291;
18516: waveform_sig_loopback =-7394;
18517: waveform_sig_loopback =-7316;
18518: waveform_sig_loopback =-6233;
18519: waveform_sig_loopback =-8217;
18520: waveform_sig_loopback =-6988;
18521: waveform_sig_loopback =-6621;
18522: waveform_sig_loopback =-7290;
18523: waveform_sig_loopback =-7804;
18524: waveform_sig_loopback =-6578;
18525: waveform_sig_loopback =-6420;
18526: waveform_sig_loopback =-8717;
18527: waveform_sig_loopback =-6364;
18528: waveform_sig_loopback =-6040;
18529: waveform_sig_loopback =-8591;
18530: waveform_sig_loopback =-7226;
18531: waveform_sig_loopback =-5672;
18532: waveform_sig_loopback =-7430;
18533: waveform_sig_loopback =-8390;
18534: waveform_sig_loopback =-5923;
18535: waveform_sig_loopback =-6542;
18536: waveform_sig_loopback =-7911;
18537: waveform_sig_loopback =-5105;
18538: waveform_sig_loopback =-10038;
18539: waveform_sig_loopback =-6838;
18540: waveform_sig_loopback =-4666;
18541: waveform_sig_loopback =-7520;
18542: waveform_sig_loopback =-7809;
18543: waveform_sig_loopback =-7929;
18544: waveform_sig_loopback =-5529;
18545: waveform_sig_loopback =-5922;
18546: waveform_sig_loopback =-8390;
18547: waveform_sig_loopback =-6695;
18548: waveform_sig_loopback =-6614;
18549: waveform_sig_loopback =-6951;
18550: waveform_sig_loopback =-6282;
18551: waveform_sig_loopback =-8230;
18552: waveform_sig_loopback =-5511;
18553: waveform_sig_loopback =-6963;
18554: waveform_sig_loopback =-7508;
18555: waveform_sig_loopback =-6095;
18556: waveform_sig_loopback =-7066;
18557: waveform_sig_loopback =-6747;
18558: waveform_sig_loopback =-7058;
18559: waveform_sig_loopback =-5685;
18560: waveform_sig_loopback =-7507;
18561: waveform_sig_loopback =-6804;
18562: waveform_sig_loopback =-5937;
18563: waveform_sig_loopback =-6759;
18564: waveform_sig_loopback =-7425;
18565: waveform_sig_loopback =-5668;
18566: waveform_sig_loopback =-6277;
18567: waveform_sig_loopback =-8007;
18568: waveform_sig_loopback =-5575;
18569: waveform_sig_loopback =-5812;
18570: waveform_sig_loopback =-7815;
18571: waveform_sig_loopback =-6530;
18572: waveform_sig_loopback =-5202;
18573: waveform_sig_loopback =-6920;
18574: waveform_sig_loopback =-7554;
18575: waveform_sig_loopback =-5230;
18576: waveform_sig_loopback =-6001;
18577: waveform_sig_loopback =-7416;
18578: waveform_sig_loopback =-4348;
18579: waveform_sig_loopback =-9180;
18580: waveform_sig_loopback =-6274;
18581: waveform_sig_loopback =-3974;
18582: waveform_sig_loopback =-6738;
18583: waveform_sig_loopback =-7191;
18584: waveform_sig_loopback =-6958;
18585: waveform_sig_loopback =-4999;
18586: waveform_sig_loopback =-5163;
18587: waveform_sig_loopback =-7404;
18588: waveform_sig_loopback =-6227;
18589: waveform_sig_loopback =-5713;
18590: waveform_sig_loopback =-6014;
18591: waveform_sig_loopback =-5720;
18592: waveform_sig_loopback =-7118;
18593: waveform_sig_loopback =-4835;
18594: waveform_sig_loopback =-6124;
18595: waveform_sig_loopback =-6342;
18596: waveform_sig_loopback =-5555;
18597: waveform_sig_loopback =-6018;
18598: waveform_sig_loopback =-5719;
18599: waveform_sig_loopback =-6380;
18600: waveform_sig_loopback =-4577;
18601: waveform_sig_loopback =-6793;
18602: waveform_sig_loopback =-5826;
18603: waveform_sig_loopback =-4714;
18604: waveform_sig_loopback =-6265;
18605: waveform_sig_loopback =-6246;
18606: waveform_sig_loopback =-4567;
18607: waveform_sig_loopback =-5588;
18608: waveform_sig_loopback =-6769;
18609: waveform_sig_loopback =-4615;
18610: waveform_sig_loopback =-4862;
18611: waveform_sig_loopback =-6706;
18612: waveform_sig_loopback =-5553;
18613: waveform_sig_loopback =-4106;
18614: waveform_sig_loopback =-5694;
18615: waveform_sig_loopback =-6777;
18616: waveform_sig_loopback =-4025;
18617: waveform_sig_loopback =-4816;
18618: waveform_sig_loopback =-6295;
18619: waveform_sig_loopback =-3218;
18620: waveform_sig_loopback =-8381;
18621: waveform_sig_loopback =-4869;
18622: waveform_sig_loopback =-2484;
18623: waveform_sig_loopback =-6090;
18624: waveform_sig_loopback =-5985;
18625: waveform_sig_loopback =-5463;
18626: waveform_sig_loopback =-4054;
18627: waveform_sig_loopback =-3693;
18628: waveform_sig_loopback =-6534;
18629: waveform_sig_loopback =-4870;
18630: waveform_sig_loopback =-4191;
18631: waveform_sig_loopback =-5190;
18632: waveform_sig_loopback =-4280;
18633: waveform_sig_loopback =-5817;
18634: waveform_sig_loopback =-3672;
18635: waveform_sig_loopback =-4809;
18636: waveform_sig_loopback =-5183;
18637: waveform_sig_loopback =-4259;
18638: waveform_sig_loopback =-4528;
18639: waveform_sig_loopback =-4653;
18640: waveform_sig_loopback =-4939;
18641: waveform_sig_loopback =-3107;
18642: waveform_sig_loopback =-5723;
18643: waveform_sig_loopback =-4300;
18644: waveform_sig_loopback =-3344;
18645: waveform_sig_loopback =-5150;
18646: waveform_sig_loopback =-4525;
18647: waveform_sig_loopback =-3348;
18648: waveform_sig_loopback =-4365;
18649: waveform_sig_loopback =-5076;
18650: waveform_sig_loopback =-3474;
18651: waveform_sig_loopback =-3308;
18652: waveform_sig_loopback =-5312;
18653: waveform_sig_loopback =-4215;
18654: waveform_sig_loopback =-2417;
18655: waveform_sig_loopback =-4499;
18656: waveform_sig_loopback =-5272;
18657: waveform_sig_loopback =-2278;
18658: waveform_sig_loopback =-3769;
18659: waveform_sig_loopback =-4544;
18660: waveform_sig_loopback =-1735;
18661: waveform_sig_loopback =-7203;
18662: waveform_sig_loopback =-2897;
18663: waveform_sig_loopback =-1229;
18664: waveform_sig_loopback =-4712;
18665: waveform_sig_loopback =-4235;
18666: waveform_sig_loopback =-4130;
18667: waveform_sig_loopback =-2420;
18668: waveform_sig_loopback =-2125;
18669: waveform_sig_loopback =-5270;
18670: waveform_sig_loopback =-3004;
18671: waveform_sig_loopback =-2763;
18672: waveform_sig_loopback =-3734;
18673: waveform_sig_loopback =-2510;
18674: waveform_sig_loopback =-4416;
18675: waveform_sig_loopback =-2012;
18676: waveform_sig_loopback =-3104;
18677: waveform_sig_loopback =-3746;
18678: waveform_sig_loopback =-2478;
18679: waveform_sig_loopback =-2913;
18680: waveform_sig_loopback =-3289;
18681: waveform_sig_loopback =-2947;
18682: waveform_sig_loopback =-1754;
18683: waveform_sig_loopback =-4143;
18684: waveform_sig_loopback =-2300;
18685: waveform_sig_loopback =-2043;
18686: waveform_sig_loopback =-3277;
18687: waveform_sig_loopback =-2895;
18688: waveform_sig_loopback =-1804;
18689: waveform_sig_loopback =-2529;
18690: waveform_sig_loopback =-3530;
18691: waveform_sig_loopback =-1696;
18692: waveform_sig_loopback =-1552;
18693: waveform_sig_loopback =-3775;
18694: waveform_sig_loopback =-2369;
18695: waveform_sig_loopback =-632;
18696: waveform_sig_loopback =-2976;
18697: waveform_sig_loopback =-3330;
18698: waveform_sig_loopback =-447;
18699: waveform_sig_loopback =-2406;
18700: waveform_sig_loopback =-2379;
18701: waveform_sig_loopback =-215;
18702: waveform_sig_loopback =-5658;
18703: waveform_sig_loopback =-522;
18704: waveform_sig_loopback =60;
18705: waveform_sig_loopback =-2760;
18706: waveform_sig_loopback =-2369;
18707: waveform_sig_loopback =-2695;
18708: waveform_sig_loopback =-47;
18709: waveform_sig_loopback =-735;
18710: waveform_sig_loopback =-3511;
18711: waveform_sig_loopback =-783;
18712: waveform_sig_loopback =-1463;
18713: waveform_sig_loopback =-1494;
18714: waveform_sig_loopback =-886;
18715: waveform_sig_loopback =-2793;
18716: waveform_sig_loopback =217;
18717: waveform_sig_loopback =-1669;
18718: waveform_sig_loopback =-1793;
18719: waveform_sig_loopback =-540;
18720: waveform_sig_loopback =-1272;
18721: waveform_sig_loopback =-1407;
18722: waveform_sig_loopback =-1037;
18723: waveform_sig_loopback =-113;
18724: waveform_sig_loopback =-2191;
18725: waveform_sig_loopback =-413;
18726: waveform_sig_loopback =-402;
18727: waveform_sig_loopback =-1278;
18728: waveform_sig_loopback =-1122;
18729: waveform_sig_loopback =69;
18730: waveform_sig_loopback =-587;
18731: waveform_sig_loopback =-1866;
18732: waveform_sig_loopback =392;
18733: waveform_sig_loopback =220;
18734: waveform_sig_loopback =-2128;
18735: waveform_sig_loopback =-156;
18736: waveform_sig_loopback =1094;
18737: waveform_sig_loopback =-1384;
18738: waveform_sig_loopback =-1213;
18739: waveform_sig_loopback =1314;
18740: waveform_sig_loopback =-598;
18741: waveform_sig_loopback =-174;
18742: waveform_sig_loopback =1169;
18743: waveform_sig_loopback =-3517;
18744: waveform_sig_loopback =1469;
18745: waveform_sig_loopback =1519;
18746: waveform_sig_loopback =-503;
18747: waveform_sig_loopback =-917;
18748: waveform_sig_loopback =-573;
18749: waveform_sig_loopback =2029;
18750: waveform_sig_loopback =622;
18751: waveform_sig_loopback =-1238;
18752: waveform_sig_loopback =928;
18753: waveform_sig_loopback =295;
18754: waveform_sig_loopback =758;
18755: waveform_sig_loopback =517;
18756: waveform_sig_loopback =-517;
18757: waveform_sig_loopback =2110;
18758: waveform_sig_loopback =-61;
18759: waveform_sig_loopback =418;
18760: waveform_sig_loopback =1080;
18761: waveform_sig_loopback =751;
18762: waveform_sig_loopback =477;
18763: waveform_sig_loopback =919;
18764: waveform_sig_loopback =1745;
18765: waveform_sig_loopback =-307;
18766: waveform_sig_loopback =1585;
18767: waveform_sig_loopback =1328;
18768: waveform_sig_loopback =822;
18769: waveform_sig_loopback =540;
18770: waveform_sig_loopback =2176;
18771: waveform_sig_loopback =1290;
18772: waveform_sig_loopback =-290;
18773: waveform_sig_loopback =2816;
18774: waveform_sig_loopback =1622;
18775: waveform_sig_loopback =-210;
18776: waveform_sig_loopback =2098;
18777: waveform_sig_loopback =2434;
18778: waveform_sig_loopback =926;
18779: waveform_sig_loopback =522;
18780: waveform_sig_loopback =3062;
18781: waveform_sig_loopback =1617;
18782: waveform_sig_loopback =1346;
18783: waveform_sig_loopback =3194;
18784: waveform_sig_loopback =-1598;
18785: waveform_sig_loopback =3230;
18786: waveform_sig_loopback =3745;
18787: waveform_sig_loopback =963;
18788: waveform_sig_loopback =976;
18789: waveform_sig_loopback =1668;
18790: waveform_sig_loopback =3513;
18791: waveform_sig_loopback =2642;
18792: waveform_sig_loopback =602;
18793: waveform_sig_loopback =2730;
18794: waveform_sig_loopback =2257;
18795: waveform_sig_loopback =2487;
18796: waveform_sig_loopback =2355;
18797: waveform_sig_loopback =1431;
18798: waveform_sig_loopback =3833;
18799: waveform_sig_loopback =1720;
18800: waveform_sig_loopback =2382;
18801: waveform_sig_loopback =2883;
18802: waveform_sig_loopback =2478;
18803: waveform_sig_loopback =2448;
18804: waveform_sig_loopback =2628;
18805: waveform_sig_loopback =3577;
18806: waveform_sig_loopback =1657;
18807: waveform_sig_loopback =3045;
18808: waveform_sig_loopback =3599;
18809: waveform_sig_loopback =2298;
18810: waveform_sig_loopback =2373;
18811: waveform_sig_loopback =4351;
18812: waveform_sig_loopback =2389;
18813: waveform_sig_loopback =2135;
18814: waveform_sig_loopback =4458;
18815: waveform_sig_loopback =3146;
18816: waveform_sig_loopback =2078;
18817: waveform_sig_loopback =3510;
18818: waveform_sig_loopback =4450;
18819: waveform_sig_loopback =2648;
18820: waveform_sig_loopback =2083;
18821: waveform_sig_loopback =5279;
18822: waveform_sig_loopback =2928;
18823: waveform_sig_loopback =3302;
18824: waveform_sig_loopback =4965;
18825: waveform_sig_loopback =-171;
18826: waveform_sig_loopback =5400;
18827: waveform_sig_loopback =5295;
18828: waveform_sig_loopback =2565;
18829: waveform_sig_loopback =2867;
18830: waveform_sig_loopback =3421;
18831: waveform_sig_loopback =5249;
18832: waveform_sig_loopback =4266;
18833: waveform_sig_loopback =2305;
18834: waveform_sig_loopback =4480;
18835: waveform_sig_loopback =4059;
18836: waveform_sig_loopback =4132;
18837: waveform_sig_loopback =3919;
18838: waveform_sig_loopback =3401;
18839: waveform_sig_loopback =5292;
18840: waveform_sig_loopback =3408;
18841: waveform_sig_loopback =4213;
18842: waveform_sig_loopback =4253;
18843: waveform_sig_loopback =4488;
18844: waveform_sig_loopback =3812;
18845: waveform_sig_loopback =4211;
18846: waveform_sig_loopback =5574;
18847: waveform_sig_loopback =2777;
18848: waveform_sig_loopback =5031;
18849: waveform_sig_loopback =5080;
18850: waveform_sig_loopback =3646;
18851: waveform_sig_loopback =4563;
18852: waveform_sig_loopback =5405;
18853: waveform_sig_loopback =4038;
18854: waveform_sig_loopback =4010;
18855: waveform_sig_loopback =5774;
18856: waveform_sig_loopback =4821;
18857: waveform_sig_loopback =3446;
18858: waveform_sig_loopback =5239;
18859: waveform_sig_loopback =6105;
18860: waveform_sig_loopback =3874;
18861: waveform_sig_loopback =3792;
18862: waveform_sig_loopback =6945;
18863: waveform_sig_loopback =4189;
18864: waveform_sig_loopback =5050;
18865: waveform_sig_loopback =6384;
18866: waveform_sig_loopback =1331;
18867: waveform_sig_loopback =7100;
18868: waveform_sig_loopback =6658;
18869: waveform_sig_loopback =3972;
18870: waveform_sig_loopback =4552;
18871: waveform_sig_loopback =4834;
18872: waveform_sig_loopback =6648;
18873: waveform_sig_loopback =5882;
18874: waveform_sig_loopback =3632;
18875: waveform_sig_loopback =5992;
18876: waveform_sig_loopback =5589;
18877: waveform_sig_loopback =5298;
18878: waveform_sig_loopback =5619;
18879: waveform_sig_loopback =4763;
18880: waveform_sig_loopback =6519;
18881: waveform_sig_loopback =5256;
18882: waveform_sig_loopback =5241;
18883: waveform_sig_loopback =5751;
18884: waveform_sig_loopback =6055;
18885: waveform_sig_loopback =4781;
18886: waveform_sig_loopback =6199;
18887: waveform_sig_loopback =6360;
18888: waveform_sig_loopback =4181;
18889: waveform_sig_loopback =6843;
18890: waveform_sig_loopback =5882;
18891: waveform_sig_loopback =5257;
18892: waveform_sig_loopback =5775;
18893: waveform_sig_loopback =6711;
18894: waveform_sig_loopback =5470;
18895: waveform_sig_loopback =5144;
18896: waveform_sig_loopback =7087;
18897: waveform_sig_loopback =6066;
18898: waveform_sig_loopback =4749;
18899: waveform_sig_loopback =6390;
18900: waveform_sig_loopback =7458;
18901: waveform_sig_loopback =4921;
18902: waveform_sig_loopback =5112;
18903: waveform_sig_loopback =8358;
18904: waveform_sig_loopback =4899;
18905: waveform_sig_loopback =6772;
18906: waveform_sig_loopback =7164;
18907: waveform_sig_loopback =2305;
18908: waveform_sig_loopback =8971;
18909: waveform_sig_loopback =7172;
18910: waveform_sig_loopback =5257;
18911: waveform_sig_loopback =5776;
18912: waveform_sig_loopback =5612;
18913: waveform_sig_loopback =8197;
18914: waveform_sig_loopback =6648;
18915: waveform_sig_loopback =4531;
18916: waveform_sig_loopback =7573;
18917: waveform_sig_loopback =6028;
18918: waveform_sig_loopback =6635;
18919: waveform_sig_loopback =6646;
18920: waveform_sig_loopback =5410;
18921: waveform_sig_loopback =7944;
18922: waveform_sig_loopback =5689;
18923: waveform_sig_loopback =6375;
18924: waveform_sig_loopback =7076;
18925: waveform_sig_loopback =6570;
18926: waveform_sig_loopback =5693;
18927: waveform_sig_loopback =7374;
18928: waveform_sig_loopback =7164;
18929: waveform_sig_loopback =5265;
18930: waveform_sig_loopback =7591;
18931: waveform_sig_loopback =6661;
18932: waveform_sig_loopback =6524;
18933: waveform_sig_loopback =6451;
18934: waveform_sig_loopback =7488;
18935: waveform_sig_loopback =6524;
18936: waveform_sig_loopback =5863;
18937: waveform_sig_loopback =8055;
18938: waveform_sig_loopback =6847;
18939: waveform_sig_loopback =5362;
18940: waveform_sig_loopback =7612;
18941: waveform_sig_loopback =8048;
18942: waveform_sig_loopback =5385;
18943: waveform_sig_loopback =6453;
18944: waveform_sig_loopback =8814;
18945: waveform_sig_loopback =5566;
18946: waveform_sig_loopback =7921;
18947: waveform_sig_loopback =7256;
18948: waveform_sig_loopback =3569;
18949: waveform_sig_loopback =9606;
18950: waveform_sig_loopback =7489;
18951: waveform_sig_loopback =6443;
18952: waveform_sig_loopback =5983;
18953: waveform_sig_loopback =6536;
18954: waveform_sig_loopback =9067;
18955: waveform_sig_loopback =6787;
18956: waveform_sig_loopback =5583;
18957: waveform_sig_loopback =8045;
18958: waveform_sig_loopback =6510;
18959: waveform_sig_loopback =7729;
18960: waveform_sig_loopback =6784;
18961: waveform_sig_loopback =6217;
18962: waveform_sig_loopback =8746;
18963: waveform_sig_loopback =6069;
18964: waveform_sig_loopback =7121;
18965: waveform_sig_loopback =7443;
18966: waveform_sig_loopback =6999;
18967: waveform_sig_loopback =6762;
18968: waveform_sig_loopback =7622;
18969: waveform_sig_loopback =7349;
18970: waveform_sig_loopback =6143;
18971: waveform_sig_loopback =7954;
18972: waveform_sig_loopback =7213;
18973: waveform_sig_loopback =6852;
18974: waveform_sig_loopback =6811;
18975: waveform_sig_loopback =8308;
18976: waveform_sig_loopback =6651;
18977: waveform_sig_loopback =6130;
18978: waveform_sig_loopback =8824;
18979: waveform_sig_loopback =6987;
18980: waveform_sig_loopback =5710;
18981: waveform_sig_loopback =8295;
18982: waveform_sig_loopback =7983;
18983: waveform_sig_loopback =6050;
18984: waveform_sig_loopback =6828;
18985: waveform_sig_loopback =8766;
18986: waveform_sig_loopback =6283;
18987: waveform_sig_loopback =8062;
18988: waveform_sig_loopback =7323;
18989: waveform_sig_loopback =4131;
18990: waveform_sig_loopback =9641;
18991: waveform_sig_loopback =7993;
18992: waveform_sig_loopback =6548;
18993: waveform_sig_loopback =5977;
18994: waveform_sig_loopback =7253;
18995: waveform_sig_loopback =8988;
18996: waveform_sig_loopback =6873;
18997: waveform_sig_loopback =6008;
18998: waveform_sig_loopback =8021;
18999: waveform_sig_loopback =6782;
19000: waveform_sig_loopback =7862;
19001: waveform_sig_loopback =6619;
19002: waveform_sig_loopback =6670;
19003: waveform_sig_loopback =8665;
19004: waveform_sig_loopback =5950;
19005: waveform_sig_loopback =7574;
19006: waveform_sig_loopback =7234;
19007: waveform_sig_loopback =7109;
19008: waveform_sig_loopback =6953;
19009: waveform_sig_loopback =7408;
19010: waveform_sig_loopback =7662;
19011: waveform_sig_loopback =6119;
19012: waveform_sig_loopback =7781;
19013: waveform_sig_loopback =7554;
19014: waveform_sig_loopback =6439;
19015: waveform_sig_loopback =7023;
19016: waveform_sig_loopback =8342;
19017: waveform_sig_loopback =6231;
19018: waveform_sig_loopback =6536;
19019: waveform_sig_loopback =8642;
19020: waveform_sig_loopback =6663;
19021: waveform_sig_loopback =5887;
19022: waveform_sig_loopback =8106;
19023: waveform_sig_loopback =7748;
19024: waveform_sig_loopback =5987;
19025: waveform_sig_loopback =6524;
19026: waveform_sig_loopback =8646;
19027: waveform_sig_loopback =6130;
19028: waveform_sig_loopback =7657;
19029: waveform_sig_loopback =7199;
19030: waveform_sig_loopback =3927;
19031: waveform_sig_loopback =9318;
19032: waveform_sig_loopback =7971;
19033: waveform_sig_loopback =5827;
19034: waveform_sig_loopback =5894;
19035: waveform_sig_loopback =7220;
19036: waveform_sig_loopback =8266;
19037: waveform_sig_loopback =6921;
19038: waveform_sig_loopback =5552;
19039: waveform_sig_loopback =7600;
19040: waveform_sig_loopback =6721;
19041: waveform_sig_loopback =7208;
19042: waveform_sig_loopback =6417;
19043: waveform_sig_loopback =6543;
19044: waveform_sig_loopback =7938;
19045: waveform_sig_loopback =5848;
19046: waveform_sig_loopback =7125;
19047: waveform_sig_loopback =6681;
19048: waveform_sig_loopback =6965;
19049: waveform_sig_loopback =6250;
19050: waveform_sig_loopback =7143;
19051: waveform_sig_loopback =7239;
19052: waveform_sig_loopback =5399;
19053: waveform_sig_loopback =7469;
19054: waveform_sig_loopback =7088;
19055: waveform_sig_loopback =5649;
19056: waveform_sig_loopback =6755;
19057: waveform_sig_loopback =7708;
19058: waveform_sig_loopback =5435;
19059: waveform_sig_loopback =6317;
19060: waveform_sig_loopback =7705;
19061: waveform_sig_loopback =6089;
19062: waveform_sig_loopback =5507;
19063: waveform_sig_loopback =7167;
19064: waveform_sig_loopback =7394;
19065: waveform_sig_loopback =5228;
19066: waveform_sig_loopback =5822;
19067: waveform_sig_loopback =8397;
19068: waveform_sig_loopback =5018;
19069: waveform_sig_loopback =7295;
19070: waveform_sig_loopback =6464;
19071: waveform_sig_loopback =2959;
19072: waveform_sig_loopback =9142;
19073: waveform_sig_loopback =6964;
19074: waveform_sig_loopback =4952;
19075: waveform_sig_loopback =5525;
19076: waveform_sig_loopback =6163;
19077: waveform_sig_loopback =7695;
19078: waveform_sig_loopback =6176;
19079: waveform_sig_loopback =4558;
19080: waveform_sig_loopback =7120;
19081: waveform_sig_loopback =5835;
19082: waveform_sig_loopback =6315;
19083: waveform_sig_loopback =5731;
19084: waveform_sig_loopback =5612;
19085: waveform_sig_loopback =7033;
19086: waveform_sig_loopback =5159;
19087: waveform_sig_loopback =6056;
19088: waveform_sig_loopback =5893;
19089: waveform_sig_loopback =6159;
19090: waveform_sig_loopback =5021;
19091: waveform_sig_loopback =6501;
19092: waveform_sig_loopback =6161;
19093: waveform_sig_loopback =4316;
19094: waveform_sig_loopback =6881;
19095: waveform_sig_loopback =5757;
19096: waveform_sig_loopback =4725;
19097: waveform_sig_loopback =6126;
19098: waveform_sig_loopback =6220;
19099: waveform_sig_loopback =4715;
19100: waveform_sig_loopback =5352;
19101: waveform_sig_loopback =6450;
19102: waveform_sig_loopback =5394;
19103: waveform_sig_loopback =4107;
19104: waveform_sig_loopback =6304;
19105: waveform_sig_loopback =6467;
19106: waveform_sig_loopback =3697;
19107: waveform_sig_loopback =5207;
19108: waveform_sig_loopback =7166;
19109: waveform_sig_loopback =3687;
19110: waveform_sig_loopback =6738;
19111: waveform_sig_loopback =4775;
19112: waveform_sig_loopback =2092;
19113: waveform_sig_loopback =8298;
19114: waveform_sig_loopback =5344;
19115: waveform_sig_loopback =4083;
19116: waveform_sig_loopback =4349;
19117: waveform_sig_loopback =4849;
19118: waveform_sig_loopback =6818;
19119: waveform_sig_loopback =4621;
19120: waveform_sig_loopback =3349;
19121: waveform_sig_loopback =6128;
19122: waveform_sig_loopback =4288;
19123: waveform_sig_loopback =5274;
19124: waveform_sig_loopback =4429;
19125: waveform_sig_loopback =4216;
19126: waveform_sig_loopback =5950;
19127: waveform_sig_loopback =3788;
19128: waveform_sig_loopback =4637;
19129: waveform_sig_loopback =4805;
19130: waveform_sig_loopback =4696;
19131: waveform_sig_loopback =3632;
19132: waveform_sig_loopback =5541;
19133: waveform_sig_loopback =4258;
19134: waveform_sig_loopback =3308;
19135: waveform_sig_loopback =5636;
19136: waveform_sig_loopback =3940;
19137: waveform_sig_loopback =3898;
19138: waveform_sig_loopback =4435;
19139: waveform_sig_loopback =4876;
19140: waveform_sig_loopback =3570;
19141: waveform_sig_loopback =3541;
19142: waveform_sig_loopback =5478;
19143: waveform_sig_loopback =3776;
19144: waveform_sig_loopback =2568;
19145: waveform_sig_loopback =5286;
19146: waveform_sig_loopback =4651;
19147: waveform_sig_loopback =2334;
19148: waveform_sig_loopback =4003;
19149: waveform_sig_loopback =5396;
19150: waveform_sig_loopback =2321;
19151: waveform_sig_loopback =5397;
19152: waveform_sig_loopback =2867;
19153: waveform_sig_loopback =920;
19154: waveform_sig_loopback =6821;
19155: waveform_sig_loopback =3579;
19156: waveform_sig_loopback =2790;
19157: waveform_sig_loopback =2623;
19158: waveform_sig_loopback =3339;
19159: waveform_sig_loopback =5550;
19160: waveform_sig_loopback =2595;
19161: waveform_sig_loopback =2079;
19162: waveform_sig_loopback =4631;
19163: waveform_sig_loopback =2313;
19164: waveform_sig_loopback =4189;
19165: waveform_sig_loopback =2399;
19166: waveform_sig_loopback =2730;
19167: waveform_sig_loopback =4608;
19168: waveform_sig_loopback =1671;
19169: waveform_sig_loopback =3435;
19170: waveform_sig_loopback =3113;
19171: waveform_sig_loopback =2762;
19172: waveform_sig_loopback =2442;
19173: waveform_sig_loopback =3623;
19174: waveform_sig_loopback =2617;
19175: waveform_sig_loopback =1950;
19176: waveform_sig_loopback =3611;
19177: waveform_sig_loopback =2540;
19178: waveform_sig_loopback =2150;
19179: waveform_sig_loopback =2652;
19180: waveform_sig_loopback =3397;
19181: waveform_sig_loopback =1657;
19182: waveform_sig_loopback =1926;
19183: waveform_sig_loopback =3943;
19184: waveform_sig_loopback =1824;
19185: waveform_sig_loopback =932;
19186: waveform_sig_loopback =3843;
19187: waveform_sig_loopback =2614;
19188: waveform_sig_loopback =733;
19189: waveform_sig_loopback =2503;
19190: waveform_sig_loopback =3305;
19191: waveform_sig_loopback =906;
19192: waveform_sig_loopback =3630;
19193: waveform_sig_loopback =760;
19194: waveform_sig_loopback =-188;
19195: waveform_sig_loopback =4671;
19196: waveform_sig_loopback =1931;
19197: waveform_sig_loopback =1176;
19198: waveform_sig_loopback =430;
19199: waveform_sig_loopback =2182;
19200: waveform_sig_loopback =3441;
19201: waveform_sig_loopback =600;
19202: waveform_sig_loopback =861;
19203: waveform_sig_loopback =2329;
19204: waveform_sig_loopback =881;
19205: waveform_sig_loopback =2446;
19206: waveform_sig_loopback =214;
19207: waveform_sig_loopback =1532;
19208: waveform_sig_loopback =2381;
19209: waveform_sig_loopback =-54;
19210: waveform_sig_loopback =1909;
19211: waveform_sig_loopback =965;
19212: waveform_sig_loopback =1193;
19213: waveform_sig_loopback =604;
19214: waveform_sig_loopback =1875;
19215: waveform_sig_loopback =738;
19216: waveform_sig_loopback =187;
19217: waveform_sig_loopback =1713;
19218: waveform_sig_loopback =890;
19219: waveform_sig_loopback =266;
19220: waveform_sig_loopback =694;
19221: waveform_sig_loopback =1865;
19222: waveform_sig_loopback =-499;
19223: waveform_sig_loopback =350;
19224: waveform_sig_loopback =2225;
19225: waveform_sig_loopback =-502;
19226: waveform_sig_loopback =-401;
19227: waveform_sig_loopback =1852;
19228: waveform_sig_loopback =489;
19229: waveform_sig_loopback =-727;
19230: waveform_sig_loopback =309;
19231: waveform_sig_loopback =1642;
19232: waveform_sig_loopback =-916;
19233: waveform_sig_loopback =1476;
19234: waveform_sig_loopback =-874;
19235: waveform_sig_loopback =-2180;
19236: waveform_sig_loopback =2824;
19237: waveform_sig_loopback =258;
19238: waveform_sig_loopback =-1121;
19239: waveform_sig_loopback =-1120;
19240: waveform_sig_loopback =407;
19241: waveform_sig_loopback =1252;
19242: waveform_sig_loopback =-987;
19243: waveform_sig_loopback =-1176;
19244: waveform_sig_loopback =412;
19245: waveform_sig_loopback =-753;
19246: waveform_sig_loopback =256;
19247: waveform_sig_loopback =-1500;
19248: waveform_sig_loopback =-206;
19249: waveform_sig_loopback =213;
19250: waveform_sig_loopback =-1719;
19251: waveform_sig_loopback =-85;
19252: waveform_sig_loopback =-939;
19253: waveform_sig_loopback =-607;
19254: waveform_sig_loopback =-1348;
19255: waveform_sig_loopback =-115;
19256: waveform_sig_loopback =-1005;
19257: waveform_sig_loopback =-1748;
19258: waveform_sig_loopback =-233;
19259: waveform_sig_loopback =-821;
19260: waveform_sig_loopback =-2046;
19261: waveform_sig_loopback =-737;
19262: waveform_sig_loopback =-130;
19263: waveform_sig_loopback =-2824;
19264: waveform_sig_loopback =-843;
19265: waveform_sig_loopback =-241;
19266: waveform_sig_loopback =-2343;
19267: waveform_sig_loopback =-1904;
19268: waveform_sig_loopback =-706;
19269: waveform_sig_loopback =-726;
19270: waveform_sig_loopback =-3262;
19271: waveform_sig_loopback =-1472;
19272: waveform_sig_loopback =231;
19273: waveform_sig_loopback =-3460;
19274: waveform_sig_loopback =47;
19275: waveform_sig_loopback =-3236;
19276: waveform_sig_loopback =-3778;
19277: waveform_sig_loopback =1292;
19278: waveform_sig_loopback =-2202;
19279: waveform_sig_loopback =-2972;
19280: waveform_sig_loopback =-2645;
19281: waveform_sig_loopback =-1532;
19282: waveform_sig_loopback =-760;
19283: waveform_sig_loopback =-2841;
19284: waveform_sig_loopback =-3001;
19285: waveform_sig_loopback =-1343;
19286: waveform_sig_loopback =-2675;
19287: waveform_sig_loopback =-1817;
19288: waveform_sig_loopback =-3093;
19289: waveform_sig_loopback =-2072;
19290: waveform_sig_loopback =-1971;
19291: waveform_sig_loopback =-3236;
19292: waveform_sig_loopback =-2067;
19293: waveform_sig_loopback =-2820;
19294: waveform_sig_loopback =-2225;
19295: waveform_sig_loopback =-3659;
19296: waveform_sig_loopback =-1472;
19297: waveform_sig_loopback =-3054;
19298: waveform_sig_loopback =-3867;
19299: waveform_sig_loopback =-1441;
19300: waveform_sig_loopback =-3253;
19301: waveform_sig_loopback =-3619;
19302: waveform_sig_loopback =-2330;
19303: waveform_sig_loopback =-2546;
19304: waveform_sig_loopback =-4112;
19305: waveform_sig_loopback =-2924;
19306: waveform_sig_loopback =-2123;
19307: waveform_sig_loopback =-3875;
19308: waveform_sig_loopback =-4080;
19309: waveform_sig_loopback =-2126;
19310: waveform_sig_loopback =-2728;
19311: waveform_sig_loopback =-5058;
19312: waveform_sig_loopback =-2905;
19313: waveform_sig_loopback =-1948;
19314: waveform_sig_loopback =-5227;
19315: waveform_sig_loopback =-1330;
19316: waveform_sig_loopback =-5346;
19317: waveform_sig_loopback =-5466;
19318: waveform_sig_loopback =-385;
19319: waveform_sig_loopback =-4080;
19320: waveform_sig_loopback =-4565;
19321: waveform_sig_loopback =-4546;
19322: waveform_sig_loopback =-3350;
19323: waveform_sig_loopback =-2168;
19324: waveform_sig_loopback =-4721;
19325: waveform_sig_loopback =-4883;
19326: waveform_sig_loopback =-2857;
19327: waveform_sig_loopback =-4465;
19328: waveform_sig_loopback =-3537;
19329: waveform_sig_loopback =-4725;
19330: waveform_sig_loopback =-3984;
19331: waveform_sig_loopback =-3340;
19332: waveform_sig_loopback =-4906;
19333: waveform_sig_loopback =-4117;
19334: waveform_sig_loopback =-4015;
19335: waveform_sig_loopback =-4196;
19336: waveform_sig_loopback =-5229;
19337: waveform_sig_loopback =-2845;
19338: waveform_sig_loopback =-5306;
19339: waveform_sig_loopback =-4896;
19340: waveform_sig_loopback =-3269;
19341: waveform_sig_loopback =-5129;
19342: waveform_sig_loopback =-4822;
19343: waveform_sig_loopback =-4325;
19344: waveform_sig_loopback =-3959;
19345: waveform_sig_loopback =-5690;
19346: waveform_sig_loopback =-4681;
19347: waveform_sig_loopback =-3436;
19348: waveform_sig_loopback =-5694;
19349: waveform_sig_loopback =-5663;
19350: waveform_sig_loopback =-3455;
19351: waveform_sig_loopback =-4497;
19352: waveform_sig_loopback =-6638;
19353: waveform_sig_loopback =-4216;
19354: waveform_sig_loopback =-3667;
19355: waveform_sig_loopback =-6717;
19356: waveform_sig_loopback =-2641;
19357: waveform_sig_loopback =-7333;
19358: waveform_sig_loopback =-6535;
19359: waveform_sig_loopback =-1829;
19360: waveform_sig_loopback =-5968;
19361: waveform_sig_loopback =-5695;
19362: waveform_sig_loopback =-6184;
19363: waveform_sig_loopback =-4795;
19364: waveform_sig_loopback =-3377;
19365: waveform_sig_loopback =-6745;
19366: waveform_sig_loopback =-5883;
19367: waveform_sig_loopback =-4279;
19368: waveform_sig_loopback =-6249;
19369: waveform_sig_loopback =-4447;
19370: waveform_sig_loopback =-6524;
19371: waveform_sig_loopback =-5266;
19372: waveform_sig_loopback =-4500;
19373: waveform_sig_loopback =-6784;
19374: waveform_sig_loopback =-5087;
19375: waveform_sig_loopback =-5456;
19376: waveform_sig_loopback =-5874;
19377: waveform_sig_loopback =-6094;
19378: waveform_sig_loopback =-4576;
19379: waveform_sig_loopback =-6544;
19380: waveform_sig_loopback =-6017;
19381: waveform_sig_loopback =-4976;
19382: waveform_sig_loopback =-6141;
19383: waveform_sig_loopback =-6239;
19384: waveform_sig_loopback =-5597;
19385: waveform_sig_loopback =-5173;
19386: waveform_sig_loopback =-7089;
19387: waveform_sig_loopback =-5912;
19388: waveform_sig_loopback =-4605;
19389: waveform_sig_loopback =-7072;
19390: waveform_sig_loopback =-6865;
19391: waveform_sig_loopback =-4429;
19392: waveform_sig_loopback =-6112;
19393: waveform_sig_loopback =-7709;
19394: waveform_sig_loopback =-5159;
19395: waveform_sig_loopback =-5332;
19396: waveform_sig_loopback =-7434;
19397: waveform_sig_loopback =-4024;
19398: waveform_sig_loopback =-8805;
19399: waveform_sig_loopback =-7042;
19400: waveform_sig_loopback =-3495;
19401: waveform_sig_loopback =-6917;
19402: waveform_sig_loopback =-6757;
19403: waveform_sig_loopback =-7691;
19404: waveform_sig_loopback =-5320;
19405: waveform_sig_loopback =-4817;
19406: waveform_sig_loopback =-7963;
19407: waveform_sig_loopback =-6512;
19408: waveform_sig_loopback =-5867;
19409: waveform_sig_loopback =-6941;
19410: waveform_sig_loopback =-5482;
19411: waveform_sig_loopback =-7932;
19412: waveform_sig_loopback =-5740;
19413: waveform_sig_loopback =-5898;
19414: waveform_sig_loopback =-7745;
19415: waveform_sig_loopback =-5841;
19416: waveform_sig_loopback =-6790;
19417: waveform_sig_loopback =-6695;
19418: waveform_sig_loopback =-6984;
19419: waveform_sig_loopback =-5757;
19420: waveform_sig_loopback =-7385;
19421: waveform_sig_loopback =-6921;
19422: waveform_sig_loopback =-6050;
19423: waveform_sig_loopback =-6873;
19424: waveform_sig_loopback =-7359;
19425: waveform_sig_loopback =-6418;
19426: waveform_sig_loopback =-5898;
19427: waveform_sig_loopback =-8294;
19428: waveform_sig_loopback =-6482;
19429: waveform_sig_loopback =-5505;
19430: waveform_sig_loopback =-8182;
19431: waveform_sig_loopback =-7333;
19432: waveform_sig_loopback =-5445;
19433: waveform_sig_loopback =-7027;
19434: waveform_sig_loopback =-8226;
19435: waveform_sig_loopback =-6144;
19436: waveform_sig_loopback =-6112;
19437: waveform_sig_loopback =-7992;
19438: waveform_sig_loopback =-5056;
19439: waveform_sig_loopback =-9454;
19440: waveform_sig_loopback =-7592;
19441: waveform_sig_loopback =-4461;
19442: waveform_sig_loopback =-7295;
19443: waveform_sig_loopback =-7870;
19444: waveform_sig_loopback =-8180;
19445: waveform_sig_loopback =-5702;
19446: waveform_sig_loopback =-6000;
19447: waveform_sig_loopback =-8265;
19448: waveform_sig_loopback =-7225;
19449: waveform_sig_loopback =-6711;
19450: waveform_sig_loopback =-7185;
19451: waveform_sig_loopback =-6548;
19452: waveform_sig_loopback =-8347;
19453: waveform_sig_loopback =-6124;
19454: waveform_sig_loopback =-6988;
19455: waveform_sig_loopback =-7910;
19456: waveform_sig_loopback =-6533;
19457: waveform_sig_loopback =-7448;
19458: waveform_sig_loopback =-6989;
19459: waveform_sig_loopback =-7701;
19460: waveform_sig_loopback =-6144;
19461: waveform_sig_loopback =-7877;
19462: waveform_sig_loopback =-7517;
19463: waveform_sig_loopback =-6375;
19464: waveform_sig_loopback =-7291;
19465: waveform_sig_loopback =-7986;
19466: waveform_sig_loopback =-6561;
19467: waveform_sig_loopback =-6523;
19468: waveform_sig_loopback =-8797;
19469: waveform_sig_loopback =-6454;
19470: waveform_sig_loopback =-6228;
19471: waveform_sig_loopback =-8559;
19472: waveform_sig_loopback =-7403;
19473: waveform_sig_loopback =-6072;
19474: waveform_sig_loopback =-7236;
19475: waveform_sig_loopback =-8559;
19476: waveform_sig_loopback =-6566;
19477: waveform_sig_loopback =-6169;
19478: waveform_sig_loopback =-8512;
19479: waveform_sig_loopback =-5300;
19480: waveform_sig_loopback =-9610;
19481: waveform_sig_loopback =-8025;
19482: waveform_sig_loopback =-4448;
19483: waveform_sig_loopback =-7646;
19484: waveform_sig_loopback =-8373;
19485: waveform_sig_loopback =-7864;
19486: waveform_sig_loopback =-6265;
19487: waveform_sig_loopback =-6118;
19488: waveform_sig_loopback =-8254;
19489: waveform_sig_loopback =-7721;
19490: waveform_sig_loopback =-6511;
19491: waveform_sig_loopback =-7411;
19492: waveform_sig_loopback =-6862;
19493: waveform_sig_loopback =-8145;
19494: waveform_sig_loopback =-6479;
19495: waveform_sig_loopback =-7059;
19496: waveform_sig_loopback =-7836;
19497: waveform_sig_loopback =-6815;
19498: waveform_sig_loopback =-7317;
19499: waveform_sig_loopback =-7083;
19500: waveform_sig_loopback =-7805;
19501: waveform_sig_loopback =-6018;
19502: waveform_sig_loopback =-7974;
19503: waveform_sig_loopback =-7572;
19504: waveform_sig_loopback =-6161;
19505: waveform_sig_loopback =-7468;
19506: waveform_sig_loopback =-7972;
19507: waveform_sig_loopback =-6187;
19508: waveform_sig_loopback =-6910;
19509: waveform_sig_loopback =-8487;
19510: waveform_sig_loopback =-6295;
19511: waveform_sig_loopback =-6500;
19512: waveform_sig_loopback =-8089;
19513: waveform_sig_loopback =-7467;
19514: waveform_sig_loopback =-5968;
19515: waveform_sig_loopback =-6878;
19516: waveform_sig_loopback =-8754;
19517: waveform_sig_loopback =-6040;
19518: waveform_sig_loopback =-6052;
19519: waveform_sig_loopback =-8586;
19520: waveform_sig_loopback =-4644;
19521: waveform_sig_loopback =-9865;
19522: waveform_sig_loopback =-7606;
19523: waveform_sig_loopback =-3905;
19524: waveform_sig_loopback =-7998;
19525: waveform_sig_loopback =-7765;
19526: waveform_sig_loopback =-7533;
19527: waveform_sig_loopback =-6289;
19528: waveform_sig_loopback =-5365;
19529: waveform_sig_loopback =-8399;
19530: waveform_sig_loopback =-7185;
19531: waveform_sig_loopback =-6017;
19532: waveform_sig_loopback =-7434;
19533: waveform_sig_loopback =-6193;
19534: waveform_sig_loopback =-7909;
19535: waveform_sig_loopback =-6073;
19536: waveform_sig_loopback =-6574;
19537: waveform_sig_loopback =-7543;
19538: waveform_sig_loopback =-6354;
19539: waveform_sig_loopback =-6852;
19540: waveform_sig_loopback =-6680;
19541: waveform_sig_loopback =-7417;
19542: waveform_sig_loopback =-5344;
19543: waveform_sig_loopback =-7683;
19544: waveform_sig_loopback =-7063;
19545: waveform_sig_loopback =-5360;
19546: waveform_sig_loopback =-7496;
19547: waveform_sig_loopback =-6983;
19548: waveform_sig_loopback =-5689;
19549: waveform_sig_loopback =-6761;
19550: waveform_sig_loopback =-7297;
19551: waveform_sig_loopback =-6234;
19552: waveform_sig_loopback =-5618;
19553: waveform_sig_loopback =-7443;
19554: waveform_sig_loopback =-7231;
19555: waveform_sig_loopback =-4662;
19556: waveform_sig_loopback =-6847;
19557: waveform_sig_loopback =-7976;
19558: waveform_sig_loopback =-4953;
19559: waveform_sig_loopback =-6086;
19560: waveform_sig_loopback =-7397;
19561: waveform_sig_loopback =-4128;
19562: waveform_sig_loopback =-9459;
19563: waveform_sig_loopback =-6265;
19564: waveform_sig_loopback =-3645;
19565: waveform_sig_loopback =-7147;
19566: waveform_sig_loopback =-6887;
19567: waveform_sig_loopback =-6956;
19568: waveform_sig_loopback =-5301;
19569: waveform_sig_loopback =-4624;
19570: waveform_sig_loopback =-7815;
19571: waveform_sig_loopback =-6095;
19572: waveform_sig_loopback =-5359;
19573: waveform_sig_loopback =-6580;
19574: waveform_sig_loopback =-5214;
19575: waveform_sig_loopback =-7228;
19576: waveform_sig_loopback =-5134;
19577: waveform_sig_loopback =-5636;
19578: waveform_sig_loopback =-6680;
19579: waveform_sig_loopback =-5565;
19580: waveform_sig_loopback =-5695;
19581: waveform_sig_loopback =-6101;
19582: waveform_sig_loopback =-6195;
19583: waveform_sig_loopback =-4398;
19584: waveform_sig_loopback =-7202;
19585: waveform_sig_loopback =-5361;
19586: waveform_sig_loopback =-5028;
19587: waveform_sig_loopback =-6336;
19588: waveform_sig_loopback =-5689;
19589: waveform_sig_loopback =-5207;
19590: waveform_sig_loopback =-5174;
19591: waveform_sig_loopback =-6698;
19592: waveform_sig_loopback =-5102;
19593: waveform_sig_loopback =-4259;
19594: waveform_sig_loopback =-6983;
19595: waveform_sig_loopback =-5744;
19596: waveform_sig_loopback =-3651;
19597: waveform_sig_loopback =-6028;
19598: waveform_sig_loopback =-6552;
19599: waveform_sig_loopback =-3986;
19600: waveform_sig_loopback =-5050;
19601: waveform_sig_loopback =-5961;
19602: waveform_sig_loopback =-3289;
19603: waveform_sig_loopback =-8399;
19604: waveform_sig_loopback =-4774;
19605: waveform_sig_loopback =-2669;
19606: waveform_sig_loopback =-5916;
19607: waveform_sig_loopback =-5705;
19608: waveform_sig_loopback =-5947;
19609: waveform_sig_loopback =-3786;
19610: waveform_sig_loopback =-3540;
19611: waveform_sig_loopback =-6844;
19612: waveform_sig_loopback =-4492;
19613: waveform_sig_loopback =-4438;
19614: waveform_sig_loopback =-5279;
19615: waveform_sig_loopback =-3795;
19616: waveform_sig_loopback =-6368;
19617: waveform_sig_loopback =-3439;
19618: waveform_sig_loopback =-4749;
19619: waveform_sig_loopback =-5496;
19620: waveform_sig_loopback =-3741;
19621: waveform_sig_loopback =-4852;
19622: waveform_sig_loopback =-4913;
19623: waveform_sig_loopback =-4459;
19624: waveform_sig_loopback =-3480;
19625: waveform_sig_loopback =-5507;
19626: waveform_sig_loopback =-4238;
19627: waveform_sig_loopback =-3838;
19628: waveform_sig_loopback =-4336;
19629: waveform_sig_loopback =-4957;
19630: waveform_sig_loopback =-3556;
19631: waveform_sig_loopback =-3757;
19632: waveform_sig_loopback =-5561;
19633: waveform_sig_loopback =-3259;
19634: waveform_sig_loopback =-3310;
19635: waveform_sig_loopback =-5449;
19636: waveform_sig_loopback =-4037;
19637: waveform_sig_loopback =-2507;
19638: waveform_sig_loopback =-4595;
19639: waveform_sig_loopback =-5033;
19640: waveform_sig_loopback =-2449;
19641: waveform_sig_loopback =-3803;
19642: waveform_sig_loopback =-4304;
19643: waveform_sig_loopback =-1976;
19644: waveform_sig_loopback =-6969;
19645: waveform_sig_loopback =-2934;
19646: waveform_sig_loopback =-1611;
19647: waveform_sig_loopback =-4148;
19648: waveform_sig_loopback =-4373;
19649: waveform_sig_loopback =-4484;
19650: waveform_sig_loopback =-1847;
19651: waveform_sig_loopback =-2614;
19652: waveform_sig_loopback =-4967;
19653: waveform_sig_loopback =-2905;
19654: waveform_sig_loopback =-3266;
19655: waveform_sig_loopback =-3110;
19656: waveform_sig_loopback =-2780;
19657: waveform_sig_loopback =-4611;
19658: waveform_sig_loopback =-1554;
19659: waveform_sig_loopback =-3525;
19660: waveform_sig_loopback =-3515;
19661: waveform_sig_loopback =-2415;
19662: waveform_sig_loopback =-3275;
19663: waveform_sig_loopback =-2790;
19664: waveform_sig_loopback =-3268;
19665: waveform_sig_loopback =-1804;
19666: waveform_sig_loopback =-3807;
19667: waveform_sig_loopback =-2681;
19668: waveform_sig_loopback =-2014;
19669: waveform_sig_loopback =-3056;
19670: waveform_sig_loopback =-3213;
19671: waveform_sig_loopback =-1727;
19672: waveform_sig_loopback =-2359;
19673: waveform_sig_loopback =-3885;
19674: waveform_sig_loopback =-1419;
19675: waveform_sig_loopback =-1702;
19676: waveform_sig_loopback =-3936;
19677: waveform_sig_loopback =-2014;
19678: waveform_sig_loopback =-1091;
19679: waveform_sig_loopback =-2760;
19680: waveform_sig_loopback =-3246;
19681: waveform_sig_loopback =-1053;
19682: waveform_sig_loopback =-1706;
19683: waveform_sig_loopback =-2773;
19684: waveform_sig_loopback =-395;
19685: waveform_sig_loopback =-5073;
19686: waveform_sig_loopback =-1368;
19687: waveform_sig_loopback =524;
19688: waveform_sig_loopback =-2696;
19689: waveform_sig_loopback =-2825;
19690: waveform_sig_loopback =-2171;
19691: waveform_sig_loopback =-383;
19692: waveform_sig_loopback =-898;
19693: waveform_sig_loopback =-2957;
19694: waveform_sig_loopback =-1333;
19695: waveform_sig_loopback =-1269;
19696: waveform_sig_loopback =-1384;
19697: waveform_sig_loopback =-1276;
19698: waveform_sig_loopback =-2295;
19699: waveform_sig_loopback =-106;
19700: waveform_sig_loopback =-1725;
19701: waveform_sig_loopback =-1421;
19702: waveform_sig_loopback =-938;
19703: waveform_sig_loopback =-1096;
19704: waveform_sig_loopback =-1183;
19705: waveform_sig_loopback =-1405;
19706: waveform_sig_loopback =153;
19707: waveform_sig_loopback =-2126;
19708: waveform_sig_loopback =-786;
19709: waveform_sig_loopback =-60;
19710: waveform_sig_loopback =-1316;
19711: waveform_sig_loopback =-1324;
19712: waveform_sig_loopback =362;
19713: waveform_sig_loopback =-883;
19714: waveform_sig_loopback =-1761;
19715: waveform_sig_loopback =560;
19716: waveform_sig_loopback =-227;
19717: waveform_sig_loopback =-1652;
19718: waveform_sig_loopback =-302;
19719: waveform_sig_loopback =716;
19720: waveform_sig_loopback =-693;
19721: waveform_sig_loopback =-1713;
19722: waveform_sig_loopback =1273;
19723: waveform_sig_loopback =-75;
19724: waveform_sig_loopback =-962;
19725: waveform_sig_loopback =1892;
19726: waveform_sig_loopback =-3663;
19727: waveform_sig_loopback =893;
19728: waveform_sig_loopback =2415;
19729: waveform_sig_loopback =-1201;
19730: waveform_sig_loopback =-612;
19731: waveform_sig_loopback =-269;
19732: waveform_sig_loopback =1321;
19733: waveform_sig_loopback =1268;
19734: waveform_sig_loopback =-1368;
19735: waveform_sig_loopback =692;
19736: waveform_sig_loopback =783;
19737: waveform_sig_loopback =243;
19738: waveform_sig_loopback =814;
19739: waveform_sig_loopback =-409;
19740: waveform_sig_loopback =1631;
19741: waveform_sig_loopback =332;
19742: waveform_sig_loopback =353;
19743: waveform_sig_loopback =921;
19744: waveform_sig_loopback =930;
19745: waveform_sig_loopback =530;
19746: waveform_sig_loopback =526;
19747: waveform_sig_loopback =2231;
19748: waveform_sig_loopback =-483;
19749: waveform_sig_loopback =1301;
19750: waveform_sig_loopback =1837;
19751: waveform_sig_loopback =211;
19752: waveform_sig_loopback =1043;
19753: waveform_sig_loopback =1993;
19754: waveform_sig_loopback =915;
19755: waveform_sig_loopback =537;
19756: waveform_sig_loopback =2051;
19757: waveform_sig_loopback =1913;
19758: waveform_sig_loopback =140;
19759: waveform_sig_loopback =1436;
19760: waveform_sig_loopback =2984;
19761: waveform_sig_loopback =778;
19762: waveform_sig_loopback =328;
19763: waveform_sig_loopback =3426;
19764: waveform_sig_loopback =1278;
19765: waveform_sig_loopback =1369;
19766: waveform_sig_loopback =3569;
19767: waveform_sig_loopback =-2013;
19768: waveform_sig_loopback =3340;
19769: waveform_sig_loopback =3873;
19770: waveform_sig_loopback =734;
19771: waveform_sig_loopback =1390;
19772: waveform_sig_loopback =1394;
19773: waveform_sig_loopback =3444;
19774: waveform_sig_loopback =3022;
19775: waveform_sig_loopback =298;
19776: waveform_sig_loopback =2801;
19777: waveform_sig_loopback =2486;
19778: waveform_sig_loopback =2070;
19779: waveform_sig_loopback =2757;
19780: waveform_sig_loopback =1287;
19781: waveform_sig_loopback =3527;
19782: waveform_sig_loopback =2298;
19783: waveform_sig_loopback =1984;
19784: waveform_sig_loopback =2828;
19785: waveform_sig_loopback =2905;
19786: waveform_sig_loopback =1972;
19787: waveform_sig_loopback =2835;
19788: waveform_sig_loopback =3697;
19789: waveform_sig_loopback =1231;
19790: waveform_sig_loopback =3600;
19791: waveform_sig_loopback =3108;
19792: waveform_sig_loopback =2414;
19793: waveform_sig_loopback =2736;
19794: waveform_sig_loopback =3633;
19795: waveform_sig_loopback =3013;
19796: waveform_sig_loopback =1976;
19797: waveform_sig_loopback =4044;
19798: waveform_sig_loopback =3657;
19799: waveform_sig_loopback =1776;
19800: waveform_sig_loopback =3439;
19801: waveform_sig_loopback =4705;
19802: waveform_sig_loopback =2384;
19803: waveform_sig_loopback =2252;
19804: waveform_sig_loopback =5271;
19805: waveform_sig_loopback =2717;
19806: waveform_sig_loopback =3555;
19807: waveform_sig_loopback =4970;
19808: waveform_sig_loopback =-388;
19809: waveform_sig_loopback =5583;
19810: waveform_sig_loopback =5112;
19811: waveform_sig_loopback =2679;
19812: waveform_sig_loopback =3066;
19813: waveform_sig_loopback =2944;
19814: waveform_sig_loopback =5546;
19815: waveform_sig_loopback =4315;
19816: waveform_sig_loopback =2048;
19817: waveform_sig_loopback =4803;
19818: waveform_sig_loopback =3785;
19819: waveform_sig_loopback =4066;
19820: waveform_sig_loopback =4378;
19821: waveform_sig_loopback =2810;
19822: waveform_sig_loopback =5543;
19823: waveform_sig_loopback =3699;
19824: waveform_sig_loopback =3656;
19825: waveform_sig_loopback =4707;
19826: waveform_sig_loopback =4260;
19827: waveform_sig_loopback =3759;
19828: waveform_sig_loopback =4621;
19829: waveform_sig_loopback =4996;
19830: waveform_sig_loopback =3176;
19831: waveform_sig_loopback =5105;
19832: waveform_sig_loopback =4613;
19833: waveform_sig_loopback =4251;
19834: waveform_sig_loopback =4065;
19835: waveform_sig_loopback =5430;
19836: waveform_sig_loopback =4583;
19837: waveform_sig_loopback =3358;
19838: waveform_sig_loopback =5942;
19839: waveform_sig_loopback =5028;
19840: waveform_sig_loopback =3246;
19841: waveform_sig_loopback =5275;
19842: waveform_sig_loopback =6049;
19843: waveform_sig_loopback =3849;
19844: waveform_sig_loopback =4045;
19845: waveform_sig_loopback =6647;
19846: waveform_sig_loopback =4175;
19847: waveform_sig_loopback =5360;
19848: waveform_sig_loopback =6055;
19849: waveform_sig_loopback =1440;
19850: waveform_sig_loopback =7106;
19851: waveform_sig_loopback =6309;
19852: waveform_sig_loopback =4510;
19853: waveform_sig_loopback =4179;
19854: waveform_sig_loopback =4620;
19855: waveform_sig_loopback =7173;
19856: waveform_sig_loopback =5386;
19857: waveform_sig_loopback =3855;
19858: waveform_sig_loopback =6117;
19859: waveform_sig_loopback =5059;
19860: waveform_sig_loopback =5849;
19861: waveform_sig_loopback =5388;
19862: waveform_sig_loopback =4464;
19863: waveform_sig_loopback =7031;
19864: waveform_sig_loopback =4686;
19865: waveform_sig_loopback =5422;
19866: waveform_sig_loopback =5957;
19867: waveform_sig_loopback =5492;
19868: waveform_sig_loopback =5311;
19869: waveform_sig_loopback =5828;
19870: waveform_sig_loopback =6324;
19871: waveform_sig_loopback =4621;
19872: waveform_sig_loopback =6292;
19873: waveform_sig_loopback =6030;
19874: waveform_sig_loopback =5509;
19875: waveform_sig_loopback =5249;
19876: waveform_sig_loopback =6935;
19877: waveform_sig_loopback =5607;
19878: waveform_sig_loopback =4658;
19879: waveform_sig_loopback =7427;
19880: waveform_sig_loopback =5953;
19881: waveform_sig_loopback =4600;
19882: waveform_sig_loopback =6733;
19883: waveform_sig_loopback =6917;
19884: waveform_sig_loopback =5251;
19885: waveform_sig_loopback =5255;
19886: waveform_sig_loopback =7723;
19887: waveform_sig_loopback =5539;
19888: waveform_sig_loopback =6383;
19889: waveform_sig_loopback =7120;
19890: waveform_sig_loopback =2765;
19891: waveform_sig_loopback =8233;
19892: waveform_sig_loopback =7544;
19893: waveform_sig_loopback =5481;
19894: waveform_sig_loopback =5190;
19895: waveform_sig_loopback =6100;
19896: waveform_sig_loopback =7996;
19897: waveform_sig_loopback =6420;
19898: waveform_sig_loopback =5084;
19899: waveform_sig_loopback =6975;
19900: waveform_sig_loopback =6264;
19901: waveform_sig_loopback =6916;
19902: waveform_sig_loopback =6197;
19903: waveform_sig_loopback =5783;
19904: waveform_sig_loopback =7879;
19905: waveform_sig_loopback =5670;
19906: waveform_sig_loopback =6684;
19907: waveform_sig_loopback =6652;
19908: waveform_sig_loopback =6655;
19909: waveform_sig_loopback =6313;
19910: waveform_sig_loopback =6625;
19911: waveform_sig_loopback =7515;
19912: waveform_sig_loopback =5420;
19913: waveform_sig_loopback =7172;
19914: waveform_sig_loopback =7207;
19915: waveform_sig_loopback =6123;
19916: waveform_sig_loopback =6494;
19917: waveform_sig_loopback =7862;
19918: waveform_sig_loopback =6144;
19919: waveform_sig_loopback =5933;
19920: waveform_sig_loopback =8196;
19921: waveform_sig_loopback =6679;
19922: waveform_sig_loopback =5636;
19923: waveform_sig_loopback =7434;
19924: waveform_sig_loopback =7821;
19925: waveform_sig_loopback =6049;
19926: waveform_sig_loopback =5964;
19927: waveform_sig_loopback =8639;
19928: waveform_sig_loopback =6260;
19929: waveform_sig_loopback =7131;
19930: waveform_sig_loopback =7889;
19931: waveform_sig_loopback =3478;
19932: waveform_sig_loopback =8991;
19933: waveform_sig_loopback =8455;
19934: waveform_sig_loopback =5829;
19935: waveform_sig_loopback =6054;
19936: waveform_sig_loopback =7023;
19937: waveform_sig_loopback =8317;
19938: waveform_sig_loopback =7474;
19939: waveform_sig_loopback =5528;
19940: waveform_sig_loopback =7690;
19941: waveform_sig_loopback =7178;
19942: waveform_sig_loopback =7184;
19943: waveform_sig_loopback =6999;
19944: waveform_sig_loopback =6451;
19945: waveform_sig_loopback =8270;
19946: waveform_sig_loopback =6489;
19947: waveform_sig_loopback =7102;
19948: waveform_sig_loopback =7201;
19949: waveform_sig_loopback =7401;
19950: waveform_sig_loopback =6582;
19951: waveform_sig_loopback =7437;
19952: waveform_sig_loopback =7907;
19953: waveform_sig_loopback =5797;
19954: waveform_sig_loopback =7938;
19955: waveform_sig_loopback =7617;
19956: waveform_sig_loopback =6430;
19957: waveform_sig_loopback =7080;
19958: waveform_sig_loopback =8308;
19959: waveform_sig_loopback =6395;
19960: waveform_sig_loopback =6626;
19961: waveform_sig_loopback =8402;
19962: waveform_sig_loopback =7046;
19963: waveform_sig_loopback =6103;
19964: waveform_sig_loopback =7645;
19965: waveform_sig_loopback =8363;
19966: waveform_sig_loopback =6237;
19967: waveform_sig_loopback =6101;
19968: waveform_sig_loopback =9312;
19969: waveform_sig_loopback =6234;
19970: waveform_sig_loopback =7757;
19971: waveform_sig_loopback =8000;
19972: waveform_sig_loopback =3371;
19973: waveform_sig_loopback =10044;
19974: waveform_sig_loopback =8367;
19975: waveform_sig_loopback =5856;
19976: waveform_sig_loopback =6561;
19977: waveform_sig_loopback =7038;
19978: waveform_sig_loopback =8820;
19979: waveform_sig_loopback =7420;
19980: waveform_sig_loopback =5444;
19981: waveform_sig_loopback =8297;
19982: waveform_sig_loopback =7087;
19983: waveform_sig_loopback =7226;
19984: waveform_sig_loopback =7252;
19985: waveform_sig_loopback =6492;
19986: waveform_sig_loopback =8480;
19987: waveform_sig_loopback =6427;
19988: waveform_sig_loopback =7112;
19989: waveform_sig_loopback =7484;
19990: waveform_sig_loopback =7342;
19991: waveform_sig_loopback =6495;
19992: waveform_sig_loopback =7628;
19993: waveform_sig_loopback =7883;
19994: waveform_sig_loopback =5675;
19995: waveform_sig_loopback =8063;
19996: waveform_sig_loopback =7452;
19997: waveform_sig_loopback =6315;
19998: waveform_sig_loopback =7388;
19999: waveform_sig_loopback =7831;
20000: waveform_sig_loopback =6487;
20001: waveform_sig_loopback =6686;
20002: waveform_sig_loopback =7999;
20003: waveform_sig_loopback =7296;
20004: waveform_sig_loopback =5693;
20005: waveform_sig_loopback =7656;
20006: waveform_sig_loopback =8481;
20007: waveform_sig_loopback =5478;
20008: waveform_sig_loopback =6642;
20009: waveform_sig_loopback =9021;
20010: waveform_sig_loopback =5553;
20011: waveform_sig_loopback =8178;
20012: waveform_sig_loopback =7196;
20013: waveform_sig_loopback =3576;
20014: waveform_sig_loopback =9799;
20015: waveform_sig_loopback =7540;
20016: waveform_sig_loopback =6179;
20017: waveform_sig_loopback =6064;
20018: waveform_sig_loopback =6630;
20019: waveform_sig_loopback =8766;
20020: waveform_sig_loopback =6842;
20021: waveform_sig_loopback =5284;
20022: waveform_sig_loopback =7938;
20023: waveform_sig_loopback =6534;
20024: waveform_sig_loopback =7182;
20025: waveform_sig_loopback =6694;
20026: waveform_sig_loopback =6064;
20027: waveform_sig_loopback =8219;
20028: waveform_sig_loopback =6010;
20029: waveform_sig_loopback =6655;
20030: waveform_sig_loopback =7019;
20031: waveform_sig_loopback =6929;
20032: waveform_sig_loopback =5894;
20033: waveform_sig_loopback =7555;
20034: waveform_sig_loopback =6892;
20035: waveform_sig_loopback =5378;
20036: waveform_sig_loopback =7933;
20037: waveform_sig_loopback =6345;
20038: waveform_sig_loopback =6329;
20039: waveform_sig_loopback =6538;
20040: waveform_sig_loopback =7298;
20041: waveform_sig_loopback =6296;
20042: waveform_sig_loopback =5514;
20043: waveform_sig_loopback =8012;
20044: waveform_sig_loopback =6486;
20045: waveform_sig_loopback =4834;
20046: waveform_sig_loopback =7631;
20047: waveform_sig_loopback =7308;
20048: waveform_sig_loopback =5061;
20049: waveform_sig_loopback =6169;
20050: waveform_sig_loopback =7969;
20051: waveform_sig_loopback =5248;
20052: waveform_sig_loopback =7430;
20053: waveform_sig_loopback =6279;
20054: waveform_sig_loopback =3132;
20055: waveform_sig_loopback =9037;
20056: waveform_sig_loopback =6842;
20057: waveform_sig_loopback =5404;
20058: waveform_sig_loopback =5277;
20059: waveform_sig_loopback =5972;
20060: waveform_sig_loopback =8091;
20061: waveform_sig_loopback =5898;
20062: waveform_sig_loopback =4556;
20063: waveform_sig_loopback =7366;
20064: waveform_sig_loopback =5376;
20065: waveform_sig_loopback =6696;
20066: waveform_sig_loopback =5712;
20067: waveform_sig_loopback =5133;
20068: waveform_sig_loopback =7692;
20069: waveform_sig_loopback =4663;
20070: waveform_sig_loopback =6046;
20071: waveform_sig_loopback =6295;
20072: waveform_sig_loopback =5539;
20073: waveform_sig_loopback =5543;
20074: waveform_sig_loopback =6394;
20075: waveform_sig_loopback =5800;
20076: waveform_sig_loopback =4935;
20077: waveform_sig_loopback =6361;
20078: waveform_sig_loopback =5815;
20079: waveform_sig_loopback =5184;
20080: waveform_sig_loopback =5368;
20081: waveform_sig_loopback =6771;
20082: waveform_sig_loopback =4725;
20083: waveform_sig_loopback =4810;
20084: waveform_sig_loopback =7098;
20085: waveform_sig_loopback =5031;
20086: waveform_sig_loopback =4037;
20087: waveform_sig_loopback =6594;
20088: waveform_sig_loopback =6065;
20089: waveform_sig_loopback =4050;
20090: waveform_sig_loopback =5119;
20091: waveform_sig_loopback =6789;
20092: waveform_sig_loopback =4191;
20093: waveform_sig_loopback =6355;
20094: waveform_sig_loopback =4841;
20095: waveform_sig_loopback =2309;
20096: waveform_sig_loopback =7839;
20097: waveform_sig_loopback =5557;
20098: waveform_sig_loopback =4309;
20099: waveform_sig_loopback =3862;
20100: waveform_sig_loopback =5140;
20101: waveform_sig_loopback =6822;
20102: waveform_sig_loopback =4327;
20103: waveform_sig_loopback =3859;
20104: waveform_sig_loopback =5822;
20105: waveform_sig_loopback =4195;
20106: waveform_sig_loopback =5732;
20107: waveform_sig_loopback =3902;
20108: waveform_sig_loopback =4528;
20109: waveform_sig_loopback =6131;
20110: waveform_sig_loopback =3224;
20111: waveform_sig_loopback =5353;
20112: waveform_sig_loopback =4457;
20113: waveform_sig_loopback =4552;
20114: waveform_sig_loopback =4257;
20115: waveform_sig_loopback =4790;
20116: waveform_sig_loopback =4870;
20117: waveform_sig_loopback =3270;
20118: waveform_sig_loopback =5126;
20119: waveform_sig_loopback =4660;
20120: waveform_sig_loopback =3443;
20121: waveform_sig_loopback =4372;
20122: waveform_sig_loopback =5244;
20123: waveform_sig_loopback =3193;
20124: waveform_sig_loopback =3662;
20125: waveform_sig_loopback =5570;
20126: waveform_sig_loopback =3538;
20127: waveform_sig_loopback =2738;
20128: waveform_sig_loopback =5226;
20129: waveform_sig_loopback =4436;
20130: waveform_sig_loopback =2778;
20131: waveform_sig_loopback =3650;
20132: waveform_sig_loopback =5294;
20133: waveform_sig_loopback =2847;
20134: waveform_sig_loopback =4693;
20135: waveform_sig_loopback =3430;
20136: waveform_sig_loopback =939;
20137: waveform_sig_loopback =6144;
20138: waveform_sig_loopback =4365;
20139: waveform_sig_loopback =2455;
20140: waveform_sig_loopback =2422;
20141: waveform_sig_loopback =3906;
20142: waveform_sig_loopback =4813;
20143: waveform_sig_loopback =3141;
20144: waveform_sig_loopback =2173;
20145: waveform_sig_loopback =4018;
20146: waveform_sig_loopback =3093;
20147: waveform_sig_loopback =3704;
20148: waveform_sig_loopback =2478;
20149: waveform_sig_loopback =3135;
20150: waveform_sig_loopback =4060;
20151: waveform_sig_loopback =2089;
20152: waveform_sig_loopback =3451;
20153: waveform_sig_loopback =2775;
20154: waveform_sig_loopback =3231;
20155: waveform_sig_loopback =2235;
20156: waveform_sig_loopback =3482;
20157: waveform_sig_loopback =3071;
20158: waveform_sig_loopback =1599;
20159: waveform_sig_loopback =3642;
20160: waveform_sig_loopback =2873;
20161: waveform_sig_loopback =1766;
20162: waveform_sig_loopback =2814;
20163: waveform_sig_loopback =3577;
20164: waveform_sig_loopback =1284;
20165: waveform_sig_loopback =2359;
20166: waveform_sig_loopback =3687;
20167: waveform_sig_loopback =1725;
20168: waveform_sig_loopback =1421;
20169: waveform_sig_loopback =3152;
20170: waveform_sig_loopback =2986;
20171: waveform_sig_loopback =949;
20172: waveform_sig_loopback =1765;
20173: waveform_sig_loopback =4016;
20174: waveform_sig_loopback =579;
20175: waveform_sig_loopback =3293;
20176: waveform_sig_loopback =1565;
20177: waveform_sig_loopback =-1073;
20178: waveform_sig_loopback =4962;
20179: waveform_sig_loopback =2205;
20180: waveform_sig_loopback =543;
20181: waveform_sig_loopback =1077;
20182: waveform_sig_loopback =1832;
20183: waveform_sig_loopback =3164;
20184: waveform_sig_loopback =1370;
20185: waveform_sig_loopback =200;
20186: waveform_sig_loopback =2550;
20187: waveform_sig_loopback =1128;
20188: waveform_sig_loopback =1813;
20189: waveform_sig_loopback =924;
20190: waveform_sig_loopback =1199;
20191: waveform_sig_loopback =2165;
20192: waveform_sig_loopback =501;
20193: waveform_sig_loopback =1377;
20194: waveform_sig_loopback =1137;
20195: waveform_sig_loopback =1429;
20196: waveform_sig_loopback =180;
20197: waveform_sig_loopback =1984;
20198: waveform_sig_loopback =983;
20199: waveform_sig_loopback =-257;
20200: waveform_sig_loopback =2066;
20201: waveform_sig_loopback =732;
20202: waveform_sig_loopback =-1;
20203: waveform_sig_loopback =1213;
20204: waveform_sig_loopback =1337;
20205: waveform_sig_loopback =-357;
20206: waveform_sig_loopback =564;
20207: waveform_sig_loopback =1590;
20208: waveform_sig_loopback =141;
20209: waveform_sig_loopback =-648;
20210: waveform_sig_loopback =1421;
20211: waveform_sig_loopback =1212;
20212: waveform_sig_loopback =-1312;
20213: waveform_sig_loopback =355;
20214: waveform_sig_loopback =2058;
20215: waveform_sig_loopback =-1562;
20216: waveform_sig_loopback =1941;
20217: waveform_sig_loopback =-799;
20218: waveform_sig_loopback =-2700;
20219: waveform_sig_loopback =3375;
20220: waveform_sig_loopback =-181;
20221: waveform_sig_loopback =-955;
20222: waveform_sig_loopback =-887;
20223: waveform_sig_loopback =-160;
20224: waveform_sig_loopback =1670;
20225: waveform_sig_loopback =-961;
20226: waveform_sig_loopback =-1527;
20227: waveform_sig_loopback =835;
20228: waveform_sig_loopback =-1021;
20229: waveform_sig_loopback =155;
20230: waveform_sig_loopback =-1080;
20231: waveform_sig_loopback =-764;
20232: waveform_sig_loopback =513;
20233: waveform_sig_loopback =-1559;
20234: waveform_sig_loopback =-550;
20235: waveform_sig_loopback =-552;
20236: waveform_sig_loopback =-669;
20237: waveform_sig_loopback =-1681;
20238: waveform_sig_loopback =353;
20239: waveform_sig_loopback =-1333;
20240: waveform_sig_loopback =-1823;
20241: waveform_sig_loopback =168;
20242: waveform_sig_loopback =-1464;
20243: waveform_sig_loopback =-1485;
20244: waveform_sig_loopback =-1000;
20245: waveform_sig_loopback =-477;
20246: waveform_sig_loopback =-2075;
20247: waveform_sig_loopback =-1672;
20248: waveform_sig_loopback =40;
20249: waveform_sig_loopback =-1968;
20250: waveform_sig_loopback =-2602;
20251: waveform_sig_loopback =-162;
20252: waveform_sig_loopback =-931;
20253: waveform_sig_loopback =-3202;
20254: waveform_sig_loopback =-1273;
20255: waveform_sig_loopback =-154;
20256: waveform_sig_loopback =-3291;
20257: waveform_sig_loopback =269;
20258: waveform_sig_loopback =-3280;
20259: waveform_sig_loopback =-4033;
20260: waveform_sig_loopback =1470;
20261: waveform_sig_loopback =-2328;
20262: waveform_sig_loopback =-2531;
20263: waveform_sig_loopback =-3057;
20264: waveform_sig_loopback =-1758;
20265: waveform_sig_loopback =-19;
20266: waveform_sig_loopback =-3325;
20267: waveform_sig_loopback =-2983;
20268: waveform_sig_loopback =-1133;
20269: waveform_sig_loopback =-2991;
20270: waveform_sig_loopback =-1378;
20271: waveform_sig_loopback =-3321;
20272: waveform_sig_loopback =-2342;
20273: waveform_sig_loopback =-1228;
20274: waveform_sig_loopback =-3726;
20275: waveform_sig_loopback =-2078;
20276: waveform_sig_loopback =-2430;
20277: waveform_sig_loopback =-2655;
20278: waveform_sig_loopback =-3228;
20279: waveform_sig_loopback =-1660;
20280: waveform_sig_loopback =-3197;
20281: waveform_sig_loopback =-3345;
20282: waveform_sig_loopback =-1938;
20283: waveform_sig_loopback =-3117;
20284: waveform_sig_loopback =-3225;
20285: waveform_sig_loopback =-2936;
20286: waveform_sig_loopback =-2059;
20287: waveform_sig_loopback =-4050;
20288: waveform_sig_loopback =-3426;
20289: waveform_sig_loopback =-1532;
20290: waveform_sig_loopback =-4083;
20291: waveform_sig_loopback =-4250;
20292: waveform_sig_loopback =-1762;
20293: waveform_sig_loopback =-3117;
20294: waveform_sig_loopback =-4699;
20295: waveform_sig_loopback =-2969;
20296: waveform_sig_loopback =-2255;
20297: waveform_sig_loopback =-4715;
20298: waveform_sig_loopback =-1628;
20299: waveform_sig_loopback =-5231;
20300: waveform_sig_loopback =-5311;
20301: waveform_sig_loopback =-719;
20302: waveform_sig_loopback =-3808;
20303: waveform_sig_loopback =-4355;
20304: waveform_sig_loopback =-4980;
20305: waveform_sig_loopback =-3051;
20306: waveform_sig_loopback =-2147;
20307: waveform_sig_loopback =-4961;
20308: waveform_sig_loopback =-4440;
20309: waveform_sig_loopback =-3198;
20310: waveform_sig_loopback =-4451;
20311: waveform_sig_loopback =-3076;
20312: waveform_sig_loopback =-5244;
20313: waveform_sig_loopback =-3711;
20314: waveform_sig_loopback =-3277;
20315: waveform_sig_loopback =-5305;
20316: waveform_sig_loopback =-3616;
20317: waveform_sig_loopback =-4357;
20318: waveform_sig_loopback =-4375;
20319: waveform_sig_loopback =-4771;
20320: waveform_sig_loopback =-3339;
20321: waveform_sig_loopback =-4860;
20322: waveform_sig_loopback =-5097;
20323: waveform_sig_loopback =-3787;
20324: waveform_sig_loopback =-4274;
20325: waveform_sig_loopback =-5184;
20326: waveform_sig_loopback =-4592;
20327: waveform_sig_loopback =-3461;
20328: waveform_sig_loopback =-5985;
20329: waveform_sig_loopback =-4546;
20330: waveform_sig_loopback =-3394;
20331: waveform_sig_loopback =-5901;
20332: waveform_sig_loopback =-5237;
20333: waveform_sig_loopback =-3706;
20334: waveform_sig_loopback =-4659;
20335: waveform_sig_loopback =-6123;
20336: waveform_sig_loopback =-4617;
20337: waveform_sig_loopback =-3578;
20338: waveform_sig_loopback =-6467;
20339: waveform_sig_loopback =-3138;
20340: waveform_sig_loopback =-6685;
20341: waveform_sig_loopback =-6858;
20342: waveform_sig_loopback =-2217;
20343: waveform_sig_loopback =-5261;
20344: waveform_sig_loopback =-6055;
20345: waveform_sig_loopback =-6302;
20346: waveform_sig_loopback =-4398;
20347: waveform_sig_loopback =-3927;
20348: waveform_sig_loopback =-6208;
20349: waveform_sig_loopback =-5953;
20350: waveform_sig_loopback =-4744;
20351: waveform_sig_loopback =-5587;
20352: waveform_sig_loopback =-4832;
20353: waveform_sig_loopback =-6527;
20354: waveform_sig_loopback =-4945;
20355: waveform_sig_loopback =-4924;
20356: waveform_sig_loopback =-6443;
20357: waveform_sig_loopback =-5079;
20358: waveform_sig_loopback =-5813;
20359: waveform_sig_loopback =-5324;
20360: waveform_sig_loopback =-6396;
20361: waveform_sig_loopback =-4788;
20362: waveform_sig_loopback =-6011;
20363: waveform_sig_loopback =-6524;
20364: waveform_sig_loopback =-4882;
20365: waveform_sig_loopback =-5840;
20366: waveform_sig_loopback =-6726;
20367: waveform_sig_loopback =-5317;
20368: waveform_sig_loopback =-5121;
20369: waveform_sig_loopback =-7365;
20370: waveform_sig_loopback =-5478;
20371: waveform_sig_loopback =-4971;
20372: waveform_sig_loopback =-6932;
20373: waveform_sig_loopback =-6551;
20374: waveform_sig_loopback =-5093;
20375: waveform_sig_loopback =-5577;
20376: waveform_sig_loopback =-7621;
20377: waveform_sig_loopback =-5726;
20378: waveform_sig_loopback =-4713;
20379: waveform_sig_loopback =-7807;
20380: waveform_sig_loopback =-4092;
20381: waveform_sig_loopback =-8208;
20382: waveform_sig_loopback =-7828;
20383: waveform_sig_loopback =-3164;
20384: waveform_sig_loopback =-6660;
20385: waveform_sig_loopback =-7312;
20386: waveform_sig_loopback =-7117;
20387: waveform_sig_loopback =-5577;
20388: waveform_sig_loopback =-5104;
20389: waveform_sig_loopback =-7246;
20390: waveform_sig_loopback =-7206;
20391: waveform_sig_loopback =-5606;
20392: waveform_sig_loopback =-6720;
20393: waveform_sig_loopback =-6136;
20394: waveform_sig_loopback =-7215;
20395: waveform_sig_loopback =-6188;
20396: waveform_sig_loopback =-6013;
20397: waveform_sig_loopback =-7252;
20398: waveform_sig_loopback =-6430;
20399: waveform_sig_loopback =-6532;
20400: waveform_sig_loopback =-6462;
20401: waveform_sig_loopback =-7505;
20402: waveform_sig_loopback =-5347;
20403: waveform_sig_loopback =-7323;
20404: waveform_sig_loopback =-7311;
20405: waveform_sig_loopback =-5653;
20406: waveform_sig_loopback =-7049;
20407: waveform_sig_loopback =-7320;
20408: waveform_sig_loopback =-6209;
20409: waveform_sig_loopback =-6241;
20410: waveform_sig_loopback =-7966;
20411: waveform_sig_loopback =-6415;
20412: waveform_sig_loopback =-5884;
20413: waveform_sig_loopback =-7687;
20414: waveform_sig_loopback =-7444;
20415: waveform_sig_loopback =-5759;
20416: waveform_sig_loopback =-6453;
20417: waveform_sig_loopback =-8604;
20418: waveform_sig_loopback =-6241;
20419: waveform_sig_loopback =-5623;
20420: waveform_sig_loopback =-8708;
20421: waveform_sig_loopback =-4560;
20422: waveform_sig_loopback =-9332;
20423: waveform_sig_loopback =-8375;
20424: waveform_sig_loopback =-3624;
20425: waveform_sig_loopback =-7859;
20426: waveform_sig_loopback =-7818;
20427: waveform_sig_loopback =-7722;
20428: waveform_sig_loopback =-6550;
20429: waveform_sig_loopback =-5342;
20430: waveform_sig_loopback =-8368;
20431: waveform_sig_loopback =-7683;
20432: waveform_sig_loopback =-5975;
20433: waveform_sig_loopback =-7812;
20434: waveform_sig_loopback =-6365;
20435: waveform_sig_loopback =-8005;
20436: waveform_sig_loopback =-6814;
20437: waveform_sig_loopback =-6376;
20438: waveform_sig_loopback =-8100;
20439: waveform_sig_loopback =-6763;
20440: waveform_sig_loopback =-7044;
20441: waveform_sig_loopback =-7191;
20442: waveform_sig_loopback =-7816;
20443: waveform_sig_loopback =-5895;
20444: waveform_sig_loopback =-7958;
20445: waveform_sig_loopback =-7651;
20446: waveform_sig_loopback =-6069;
20447: waveform_sig_loopback =-7714;
20448: waveform_sig_loopback =-7607;
20449: waveform_sig_loopback =-6618;
20450: waveform_sig_loopback =-6874;
20451: waveform_sig_loopback =-8106;
20452: waveform_sig_loopback =-7085;
20453: waveform_sig_loopback =-6139;
20454: waveform_sig_loopback =-8040;
20455: waveform_sig_loopback =-8141;
20456: waveform_sig_loopback =-5652;
20457: waveform_sig_loopback =-7189;
20458: waveform_sig_loopback =-8935;
20459: waveform_sig_loopback =-6117;
20460: waveform_sig_loopback =-6523;
20461: waveform_sig_loopback =-8580;
20462: waveform_sig_loopback =-4879;
20463: waveform_sig_loopback =-10046;
20464: waveform_sig_loopback =-7943;
20465: waveform_sig_loopback =-4299;
20466: waveform_sig_loopback =-8014;
20467: waveform_sig_loopback =-7806;
20468: waveform_sig_loopback =-8321;
20469: waveform_sig_loopback =-6374;
20470: waveform_sig_loopback =-5600;
20471: waveform_sig_loopback =-8815;
20472: waveform_sig_loopback =-7486;
20473: waveform_sig_loopback =-6386;
20474: waveform_sig_loopback =-7846;
20475: waveform_sig_loopback =-6330;
20476: waveform_sig_loopback =-8466;
20477: waveform_sig_loopback =-6587;
20478: waveform_sig_loopback =-6566;
20479: waveform_sig_loopback =-8291;
20480: waveform_sig_loopback =-6714;
20481: waveform_sig_loopback =-7151;
20482: waveform_sig_loopback =-7302;
20483: waveform_sig_loopback =-7728;
20484: waveform_sig_loopback =-5919;
20485: waveform_sig_loopback =-8169;
20486: waveform_sig_loopback =-7303;
20487: waveform_sig_loopback =-6361;
20488: waveform_sig_loopback =-7657;
20489: waveform_sig_loopback =-7389;
20490: waveform_sig_loopback =-6945;
20491: waveform_sig_loopback =-6487;
20492: waveform_sig_loopback =-8251;
20493: waveform_sig_loopback =-7045;
20494: waveform_sig_loopback =-5692;
20495: waveform_sig_loopback =-8450;
20496: waveform_sig_loopback =-7632;
20497: waveform_sig_loopback =-5457;
20498: waveform_sig_loopback =-7415;
20499: waveform_sig_loopback =-8344;
20500: waveform_sig_loopback =-6114;
20501: waveform_sig_loopback =-6427;
20502: waveform_sig_loopback =-8014;
20503: waveform_sig_loopback =-5081;
20504: waveform_sig_loopback =-9717;
20505: waveform_sig_loopback =-7518;
20506: waveform_sig_loopback =-4319;
20507: waveform_sig_loopback =-7553;
20508: waveform_sig_loopback =-7784;
20509: waveform_sig_loopback =-7954;
20510: waveform_sig_loopback =-5939;
20511: waveform_sig_loopback =-5444;
20512: waveform_sig_loopback =-8486;
20513: waveform_sig_loopback =-7076;
20514: waveform_sig_loopback =-6193;
20515: waveform_sig_loopback =-7436;
20516: waveform_sig_loopback =-5889;
20517: waveform_sig_loopback =-8330;
20518: waveform_sig_loopback =-5936;
20519: waveform_sig_loopback =-6310;
20520: waveform_sig_loopback =-7989;
20521: waveform_sig_loopback =-5985;
20522: waveform_sig_loopback =-6961;
20523: waveform_sig_loopback =-6920;
20524: waveform_sig_loopback =-6911;
20525: waveform_sig_loopback =-5909;
20526: waveform_sig_loopback =-7441;
20527: waveform_sig_loopback =-6784;
20528: waveform_sig_loopback =-6128;
20529: waveform_sig_loopback =-6663;
20530: waveform_sig_loopback =-7379;
20531: waveform_sig_loopback =-5974;
20532: waveform_sig_loopback =-5965;
20533: waveform_sig_loopback =-8121;
20534: waveform_sig_loopback =-5813;
20535: waveform_sig_loopback =-5548;
20536: waveform_sig_loopback =-7834;
20537: waveform_sig_loopback =-6771;
20538: waveform_sig_loopback =-5077;
20539: waveform_sig_loopback =-6680;
20540: waveform_sig_loopback =-7756;
20541: waveform_sig_loopback =-5387;
20542: waveform_sig_loopback =-5794;
20543: waveform_sig_loopback =-7317;
20544: waveform_sig_loopback =-4420;
20545: waveform_sig_loopback =-9179;
20546: waveform_sig_loopback =-6499;
20547: waveform_sig_loopback =-3767;
20548: waveform_sig_loopback =-6787;
20549: waveform_sig_loopback =-7140;
20550: waveform_sig_loopback =-7156;
20551: waveform_sig_loopback =-4887;
20552: waveform_sig_loopback =-5090;
20553: waveform_sig_loopback =-7556;
20554: waveform_sig_loopback =-6010;
20555: waveform_sig_loopback =-5730;
20556: waveform_sig_loopback =-6263;
20557: waveform_sig_loopback =-5392;
20558: waveform_sig_loopback =-7353;
20559: waveform_sig_loopback =-4797;
20560: waveform_sig_loopback =-6019;
20561: waveform_sig_loopback =-6675;
20562: waveform_sig_loopback =-5167;
20563: waveform_sig_loopback =-6309;
20564: waveform_sig_loopback =-5645;
20565: waveform_sig_loopback =-6330;
20566: waveform_sig_loopback =-4808;
20567: waveform_sig_loopback =-6415;
20568: waveform_sig_loopback =-6127;
20569: waveform_sig_loopback =-4777;
20570: waveform_sig_loopback =-5972;
20571: waveform_sig_loopback =-6411;
20572: waveform_sig_loopback =-4684;
20573: waveform_sig_loopback =-5399;
20574: waveform_sig_loopback =-6883;
20575: waveform_sig_loopback =-4757;
20576: waveform_sig_loopback =-4652;
20577: waveform_sig_loopback =-6796;
20578: waveform_sig_loopback =-5653;
20579: waveform_sig_loopback =-4024;
20580: waveform_sig_loopback =-5730;
20581: waveform_sig_loopback =-6604;
20582: waveform_sig_loopback =-4385;
20583: waveform_sig_loopback =-4606;
20584: waveform_sig_loopback =-6249;
20585: waveform_sig_loopback =-3408;
20586: waveform_sig_loopback =-7873;
20587: waveform_sig_loopback =-5393;
20588: waveform_sig_loopback =-2515;
20589: waveform_sig_loopback =-5641;
20590: waveform_sig_loopback =-6229;
20591: waveform_sig_loopback =-5543;
20592: waveform_sig_loopback =-3848;
20593: waveform_sig_loopback =-3926;
20594: waveform_sig_loopback =-6144;
20595: waveform_sig_loopback =-5144;
20596: waveform_sig_loopback =-4285;
20597: waveform_sig_loopback =-4938;
20598: waveform_sig_loopback =-4479;
20599: waveform_sig_loopback =-5704;
20600: waveform_sig_loopback =-3700;
20601: waveform_sig_loopback =-4797;
20602: waveform_sig_loopback =-5067;
20603: waveform_sig_loopback =-4302;
20604: waveform_sig_loopback =-4623;
20605: waveform_sig_loopback =-4462;
20606: waveform_sig_loopback =-5111;
20607: waveform_sig_loopback =-3037;
20608: waveform_sig_loopback =-5473;
20609: waveform_sig_loopback =-4516;
20610: waveform_sig_loopback =-3407;
20611: waveform_sig_loopback =-4818;
20612: waveform_sig_loopback =-4869;
20613: waveform_sig_loopback =-3266;
20614: waveform_sig_loopback =-4096;
20615: waveform_sig_loopback =-5354;
20616: waveform_sig_loopback =-3298;
20617: waveform_sig_loopback =-3381;
20618: waveform_sig_loopback =-5240;
20619: waveform_sig_loopback =-4181;
20620: waveform_sig_loopback =-2704;
20621: waveform_sig_loopback =-4069;
20622: waveform_sig_loopback =-5327;
20623: waveform_sig_loopback =-2704;
20624: waveform_sig_loopback =-3115;
20625: waveform_sig_loopback =-5071;
20626: waveform_sig_loopback =-1530;
20627: waveform_sig_loopback =-6725;
20628: waveform_sig_loopback =-3760;
20629: waveform_sig_loopback =-649;
20630: waveform_sig_loopback =-4677;
20631: waveform_sig_loopback =-4327;
20632: waveform_sig_loopback =-3919;
20633: waveform_sig_loopback =-2722;
20634: waveform_sig_loopback =-1939;
20635: waveform_sig_loopback =-4975;
20636: waveform_sig_loopback =-3365;
20637: waveform_sig_loopback =-2519;
20638: waveform_sig_loopback =-3739;
20639: waveform_sig_loopback =-2586;
20640: waveform_sig_loopback =-4192;
20641: waveform_sig_loopback =-2242;
20642: waveform_sig_loopback =-2966;
20643: waveform_sig_loopback =-3584;
20644: waveform_sig_loopback =-2673;
20645: waveform_sig_loopback =-2825;
20646: waveform_sig_loopback =-3008;
20647: waveform_sig_loopback =-3339;
20648: waveform_sig_loopback =-1421;
20649: waveform_sig_loopback =-4040;
20650: waveform_sig_loopback =-2631;
20651: waveform_sig_loopback =-1653;
20652: waveform_sig_loopback =-3433;
20653: waveform_sig_loopback =-2846;
20654: waveform_sig_loopback =-1743;
20655: waveform_sig_loopback =-2597;
20656: waveform_sig_loopback =-3338;
20657: waveform_sig_loopback =-1845;
20658: waveform_sig_loopback =-1553;
20659: waveform_sig_loopback =-3454;
20660: waveform_sig_loopback =-2666;
20661: waveform_sig_loopback =-708;
20662: waveform_sig_loopback =-2600;
20663: waveform_sig_loopback =-3700;
20664: waveform_sig_loopback =-497;
20665: waveform_sig_loopback =-2085;
20666: waveform_sig_loopback =-2966;
20667: waveform_sig_loopback =435;
20668: waveform_sig_loopback =-5561;
20669: waveform_sig_loopback =-1482;
20670: waveform_sig_loopback =644;
20671: waveform_sig_loopback =-2856;
20672: waveform_sig_loopback =-2249;
20673: waveform_sig_loopback =-2684;
20674: waveform_sig_loopback =-690;
20675: waveform_sig_loopback =-54;
20676: waveform_sig_loopback =-3574;
20677: waveform_sig_loopback =-1320;
20678: waveform_sig_loopback =-947;
20679: waveform_sig_loopback =-1927;
20680: waveform_sig_loopback =-597;
20681: waveform_sig_loopback =-2768;
20682: waveform_sig_loopback =-252;
20683: waveform_sig_loopback =-1118;
20684: waveform_sig_loopback =-2053;
20685: waveform_sig_loopback =-753;
20686: waveform_sig_loopback =-1054;
20687: waveform_sig_loopback =-1373;
20688: waveform_sig_loopback =-1243;
20689: waveform_sig_loopback =147;
20690: waveform_sig_loopback =-2360;
20691: waveform_sig_loopback =-426;
20692: waveform_sig_loopback =-230;
20693: waveform_sig_loopback =-1513;
20694: waveform_sig_loopback =-869;
20695: waveform_sig_loopback =-107;
20696: waveform_sig_loopback =-548;
20697: waveform_sig_loopback =-1740;
20698: waveform_sig_loopback =25;
20699: waveform_sig_loopback =434;
20700: waveform_sig_loopback =-1970;
20701: waveform_sig_loopback =-634;
20702: waveform_sig_loopback =1343;
20703: waveform_sig_loopback =-1107;
20704: waveform_sig_loopback =-1585;
20705: waveform_sig_loopback =1413;
20706: waveform_sig_loopback =-458;
20707: waveform_sig_loopback =-586;
20708: waveform_sig_loopback =1735;
20709: waveform_sig_loopback =-3767;
20710: waveform_sig_loopback =1168;
20711: waveform_sig_loopback =1942;
20712: waveform_sig_loopback =-828;
20713: waveform_sig_loopback =-463;
20714: waveform_sig_loopback =-885;
20715: waveform_sig_loopback =1832;
20716: waveform_sig_loopback =1184;
20717: waveform_sig_loopback =-1600;
20718: waveform_sig_loopback =990;
20719: waveform_sig_loopback =479;
20720: waveform_sig_loopback =319;
20721: waveform_sig_loopback =1073;
20722: waveform_sig_loopback =-913;
20723: waveform_sig_loopback =2021;
20724: waveform_sig_loopback =356;
20725: waveform_sig_loopback =-5;
20726: waveform_sig_loopback =1334;
20727: waveform_sig_loopback =659;
20728: waveform_sig_loopback =504;
20729: waveform_sig_loopback =814;
20730: waveform_sig_loopback =1815;
20731: waveform_sig_loopback =-331;
20732: waveform_sig_loopback =1511;
20733: waveform_sig_loopback =1395;
20734: waveform_sig_loopback =728;
20735: waveform_sig_loopback =750;
20736: waveform_sig_loopback =1822;
20737: waveform_sig_loopback =1553;
20738: waveform_sig_loopback =-172;
20739: waveform_sig_loopback =2294;
20740: waveform_sig_loopback =2192;
20741: waveform_sig_loopback =-308;
20742: waveform_sig_loopback =1740;
20743: waveform_sig_loopback =2886;
20744: waveform_sig_loopback =711;
20745: waveform_sig_loopback =631;
20746: waveform_sig_loopback =3033;
20747: waveform_sig_loopback =1518;
20748: waveform_sig_loopback =1489;
20749: waveform_sig_loopback =3196;
20750: waveform_sig_loopback =-1591;
20751: waveform_sig_loopback =3066;
20752: waveform_sig_loopback =3620;
20753: waveform_sig_loopback =1384;
20754: waveform_sig_loopback =972;
20755: waveform_sig_loopback =1308;
20756: waveform_sig_loopback =3783;
20757: waveform_sig_loopback =2604;
20758: waveform_sig_loopback =698;
20759: waveform_sig_loopback =2640;
20760: waveform_sig_loopback =2296;
20761: waveform_sig_loopback =2484;
20762: waveform_sig_loopback =2536;
20763: waveform_sig_loopback =1196;
20764: waveform_sig_loopback =3864;
20765: waveform_sig_loopback =2034;
20766: waveform_sig_loopback =2073;
20767: waveform_sig_loopback =3036;
20768: waveform_sig_loopback =2485;
20769: waveform_sig_loopback =2386;
20770: waveform_sig_loopback =2729;
20771: waveform_sig_loopback =3458;
20772: waveform_sig_loopback =1716;
20773: waveform_sig_loopback =3204;
20774: waveform_sig_loopback =3199;
20775: waveform_sig_loopback =2777;
20776: waveform_sig_loopback =2178;
20777: waveform_sig_loopback =4054;
20778: waveform_sig_loopback =3085;
20779: waveform_sig_loopback =1463;
20780: waveform_sig_loopback =4641;
20781: waveform_sig_loopback =3350;
20782: waveform_sig_loopback =1748;
20783: waveform_sig_loopback =3705;
20784: waveform_sig_loopback =4216;
20785: waveform_sig_loopback =2892;
20786: waveform_sig_loopback =2082;
20787: waveform_sig_loopback =4869;
20788: waveform_sig_loopback =3389;
20789: waveform_sig_loopback =2963;
20790: waveform_sig_loopback =5148;
20791: waveform_sig_loopback =-22;
20792: waveform_sig_loopback =4868;
20793: waveform_sig_loopback =5545;
20794: waveform_sig_loopback =2695;
20795: waveform_sig_loopback =2802;
20796: waveform_sig_loopback =3306;
20797: waveform_sig_loopback =5241;
20798: waveform_sig_loopback =4328;
20799: waveform_sig_loopback =2403;
20800: waveform_sig_loopback =4431;
20801: waveform_sig_loopback =4044;
20802: waveform_sig_loopback =4119;
20803: waveform_sig_loopback =4086;
20804: waveform_sig_loopback =3193;
20805: waveform_sig_loopback =5480;
20806: waveform_sig_loopback =3651;
20807: waveform_sig_loopback =3877;
20808: waveform_sig_loopback =4455;
20809: waveform_sig_loopback =4195;
20810: waveform_sig_loopback =4283;
20811: waveform_sig_loopback =4106;
20812: waveform_sig_loopback =5240;
20813: waveform_sig_loopback =3166;
20814: waveform_sig_loopback =4735;
20815: waveform_sig_loopback =5349;
20816: waveform_sig_loopback =3654;
20817: waveform_sig_loopback =4020;
20818: waveform_sig_loopback =5847;
20819: waveform_sig_loopback =4156;
20820: waveform_sig_loopback =3667;
20821: waveform_sig_loopback =5689;
20822: waveform_sig_loopback =5001;
20823: waveform_sig_loopback =3541;
20824: waveform_sig_loopback =4855;
20825: waveform_sig_loopback =6168;
20826: waveform_sig_loopback =4246;
20827: waveform_sig_loopback =3527;
20828: waveform_sig_loopback =6706;
20829: waveform_sig_loopback =4608;
20830: waveform_sig_loopback =4809;
20831: waveform_sig_loopback =6618;
20832: waveform_sig_loopback =1252;
20833: waveform_sig_loopback =6824;
20834: waveform_sig_loopback =6945;
20835: waveform_sig_loopback =3938;
20836: waveform_sig_loopback =4445;
20837: waveform_sig_loopback =4817;
20838: waveform_sig_loopback =6660;
20839: waveform_sig_loopback =5876;
20840: waveform_sig_loopback =3734;
20841: waveform_sig_loopback =5854;
20842: waveform_sig_loopback =5576;
20843: waveform_sig_loopback =5307;
20844: waveform_sig_loopback =5540;
20845: waveform_sig_loopback =4727;
20846: waveform_sig_loopback =6560;
20847: waveform_sig_loopback =5125;
20848: waveform_sig_loopback =5296;
20849: waveform_sig_loopback =5713;
20850: waveform_sig_loopback =5946;
20851: waveform_sig_loopback =4950;
20852: waveform_sig_loopback =5674;
20853: waveform_sig_loopback =6905;
20854: waveform_sig_loopback =4007;
20855: waveform_sig_loopback =6471;
20856: waveform_sig_loopback =6212;
20857: waveform_sig_loopback =5133;
20858: waveform_sig_loopback =5774;
20859: waveform_sig_loopback =6506;
20860: waveform_sig_loopback =5746;
20861: waveform_sig_loopback =4988;
20862: waveform_sig_loopback =6879;
20863: waveform_sig_loopback =6404;
20864: waveform_sig_loopback =4576;
20865: waveform_sig_loopback =6369;
20866: waveform_sig_loopback =7289;
20867: waveform_sig_loopback =5184;
20868: waveform_sig_loopback =5033;
20869: waveform_sig_loopback =7959;
20870: waveform_sig_loopback =5488;
20871: waveform_sig_loopback =6163;
20872: waveform_sig_loopback =7611;
20873: waveform_sig_loopback =2360;
20874: waveform_sig_loopback =8186;
20875: waveform_sig_loopback =7848;
20876: waveform_sig_loopback =5122;
20877: waveform_sig_loopback =5635;
20878: waveform_sig_loopback =5744;
20879: waveform_sig_loopback =7857;
20880: waveform_sig_loopback =7068;
20881: waveform_sig_loopback =4443;
20882: waveform_sig_loopback =7202;
20883: waveform_sig_loopback =6493;
20884: waveform_sig_loopback =6398;
20885: waveform_sig_loopback =6813;
20886: waveform_sig_loopback =5289;
20887: waveform_sig_loopback =7878;
20888: waveform_sig_loopback =6153;
20889: waveform_sig_loopback =5962;
20890: waveform_sig_loopback =7094;
20891: waveform_sig_loopback =6664;
20892: waveform_sig_loopback =5967;
20893: waveform_sig_loopback =7023;
20894: waveform_sig_loopback =7285;
20895: waveform_sig_loopback =5396;
20896: waveform_sig_loopback =7381;
20897: waveform_sig_loopback =6919;
20898: waveform_sig_loopback =6308;
20899: waveform_sig_loopback =6406;
20900: waveform_sig_loopback =7681;
20901: waveform_sig_loopback =6478;
20902: waveform_sig_loopback =5787;
20903: waveform_sig_loopback =7930;
20904: waveform_sig_loopback =7133;
20905: waveform_sig_loopback =5414;
20906: waveform_sig_loopback =7208;
20907: waveform_sig_loopback =8225;
20908: waveform_sig_loopback =5729;
20909: waveform_sig_loopback =6047;
20910: waveform_sig_loopback =8761;
20911: waveform_sig_loopback =5906;
20912: waveform_sig_loopback =7450;
20913: waveform_sig_loopback =7866;
20914: waveform_sig_loopback =3184;
20915: waveform_sig_loopback =9304;
20916: waveform_sig_loopback =8042;
20917: waveform_sig_loopback =6131;
20918: waveform_sig_loopback =6161;
20919: waveform_sig_loopback =6364;
20920: waveform_sig_loopback =8926;
20921: waveform_sig_loopback =7114;
20922: waveform_sig_loopback =5360;
20923: waveform_sig_loopback =8016;
20924: waveform_sig_loopback =6685;
20925: waveform_sig_loopback =7391;
20926: waveform_sig_loopback =7071;
20927: waveform_sig_loopback =5963;
20928: waveform_sig_loopback =8721;
20929: waveform_sig_loopback =6278;
20930: waveform_sig_loopback =6856;
20931: waveform_sig_loopback =7584;
20932: waveform_sig_loopback =7029;
20933: waveform_sig_loopback =6695;
20934: waveform_sig_loopback =7439;
20935: waveform_sig_loopback =7695;
20936: waveform_sig_loopback =6004;
20937: waveform_sig_loopback =7802;
20938: waveform_sig_loopback =7401;
20939: waveform_sig_loopback =6798;
20940: waveform_sig_loopback =6785;
20941: waveform_sig_loopback =8140;
20942: waveform_sig_loopback =6895;
20943: waveform_sig_loopback =6119;
20944: waveform_sig_loopback =8515;
20945: waveform_sig_loopback =7366;
20946: waveform_sig_loopback =5675;
20947: waveform_sig_loopback =7940;
20948: waveform_sig_loopback =8287;
20949: waveform_sig_loopback =6014;
20950: waveform_sig_loopback =6711;
20951: waveform_sig_loopback =8783;
20952: waveform_sig_loopback =6360;
20953: waveform_sig_loopback =7847;
20954: waveform_sig_loopback =7741;
20955: waveform_sig_loopback =3937;
20956: waveform_sig_loopback =9342;
20957: waveform_sig_loopback =8323;
20958: waveform_sig_loopback =6571;
20959: waveform_sig_loopback =5991;
20960: waveform_sig_loopback =7001;
20961: waveform_sig_loopback =9093;
20962: waveform_sig_loopback =7185;
20963: waveform_sig_loopback =5820;
20964: waveform_sig_loopback =7960;
20965: waveform_sig_loopback =6971;
20966: waveform_sig_loopback =7783;
20967: waveform_sig_loopback =6898;
20968: waveform_sig_loopback =6406;
20969: waveform_sig_loopback =8803;
20970: waveform_sig_loopback =6263;
20971: waveform_sig_loopback =7266;
20972: waveform_sig_loopback =7461;
20973: waveform_sig_loopback =7160;
20974: waveform_sig_loopback =6875;
20975: waveform_sig_loopback =7463;
20976: waveform_sig_loopback =7697;
20977: waveform_sig_loopback =6146;
20978: waveform_sig_loopback =7731;
20979: waveform_sig_loopback =7513;
20980: waveform_sig_loopback =6688;
20981: waveform_sig_loopback =6687;
20982: waveform_sig_loopback =8442;
20983: waveform_sig_loopback =6474;
20984: waveform_sig_loopback =6146;
20985: waveform_sig_loopback =8692;
20986: waveform_sig_loopback =6882;
20987: waveform_sig_loopback =5876;
20988: waveform_sig_loopback =7814;
20989: waveform_sig_loopback =7986;
20990: waveform_sig_loopback =6142;
20991: waveform_sig_loopback =6352;
20992: waveform_sig_loopback =8736;
20993: waveform_sig_loopback =6246;
20994: waveform_sig_loopback =7580;
20995: waveform_sig_loopback =7577;
20996: waveform_sig_loopback =3702;
20997: waveform_sig_loopback =9234;
20998: waveform_sig_loopback =8159;
20999: waveform_sig_loopback =6000;
21000: waveform_sig_loopback =5884;
21001: waveform_sig_loopback =6978;
21002: waveform_sig_loopback =8471;
21003: waveform_sig_loopback =6975;
21004: waveform_sig_loopback =5526;
21005: waveform_sig_loopback =7655;
21006: waveform_sig_loopback =6674;
21007: waveform_sig_loopback =7343;
21008: waveform_sig_loopback =6473;
21009: waveform_sig_loopback =6205;
21010: waveform_sig_loopback =8269;
21011: waveform_sig_loopback =5715;
21012: waveform_sig_loopback =7114;
21013: waveform_sig_loopback =6683;
21014: waveform_sig_loopback =6771;
21015: waveform_sig_loopback =6530;
21016: waveform_sig_loopback =6829;
21017: waveform_sig_loopback =7444;
21018: waveform_sig_loopback =5215;
21019: waveform_sig_loopback =7500;
21020: waveform_sig_loopback =7245;
21021: waveform_sig_loopback =5693;
21022: waveform_sig_loopback =6459;
21023: waveform_sig_loopback =7766;
21024: waveform_sig_loopback =5892;
21025: waveform_sig_loopback =5794;
21026: waveform_sig_loopback =7788;
21027: waveform_sig_loopback =6411;
21028: waveform_sig_loopback =5338;
21029: waveform_sig_loopback =7113;
21030: waveform_sig_loopback =7315;
21031: waveform_sig_loopback =5515;
21032: waveform_sig_loopback =5731;
21033: waveform_sig_loopback =8110;
21034: waveform_sig_loopback =5409;
21035: waveform_sig_loopback =6996;
21036: waveform_sig_loopback =6874;
21037: waveform_sig_loopback =2820;
21038: waveform_sig_loopback =8722;
21039: waveform_sig_loopback =7442;
21040: waveform_sig_loopback =4991;
21041: waveform_sig_loopback =5319;
21042: waveform_sig_loopback =6215;
21043: waveform_sig_loopback =7614;
21044: waveform_sig_loopback =6333;
21045: waveform_sig_loopback =4480;
21046: waveform_sig_loopback =6952;
21047: waveform_sig_loopback =5945;
21048: waveform_sig_loopback =6286;
21049: waveform_sig_loopback =5770;
21050: waveform_sig_loopback =5435;
21051: waveform_sig_loopback =7218;
21052: waveform_sig_loopback =5083;
21053: waveform_sig_loopback =6014;
21054: waveform_sig_loopback =5896;
21055: waveform_sig_loopback =6144;
21056: waveform_sig_loopback =5169;
21057: waveform_sig_loopback =6182;
21058: waveform_sig_loopback =6498;
21059: waveform_sig_loopback =4267;
21060: waveform_sig_loopback =6608;
21061: waveform_sig_loopback =6002;
21062: waveform_sig_loopback =4798;
21063: waveform_sig_loopback =5825;
21064: waveform_sig_loopback =6421;
21065: waveform_sig_loopback =4839;
21066: waveform_sig_loopback =5106;
21067: waveform_sig_loopback =6581;
21068: waveform_sig_loopback =5421;
21069: waveform_sig_loopback =4186;
21070: waveform_sig_loopback =6133;
21071: waveform_sig_loopback =6423;
21072: waveform_sig_loopback =4064;
21073: waveform_sig_loopback =4803;
21074: waveform_sig_loopback =7194;
21075: waveform_sig_loopback =3996;
21076: waveform_sig_loopback =6161;
21077: waveform_sig_loopback =5480;
21078: waveform_sig_loopback =1702;
21079: waveform_sig_loopback =7942;
21080: waveform_sig_loopback =5881;
21081: waveform_sig_loopback =3867;
21082: waveform_sig_loopback =4389;
21083: waveform_sig_loopback =4828;
21084: waveform_sig_loopback =6589;
21085: waveform_sig_loopback =4995;
21086: waveform_sig_loopback =3211;
21087: waveform_sig_loopback =6032;
21088: waveform_sig_loopback =4438;
21089: waveform_sig_loopback =5132;
21090: waveform_sig_loopback =4627;
21091: waveform_sig_loopback =4018;
21092: waveform_sig_loopback =6028;
21093: waveform_sig_loopback =3805;
21094: waveform_sig_loopback =4624;
21095: waveform_sig_loopback =4790;
21096: waveform_sig_loopback =4719;
21097: waveform_sig_loopback =3764;
21098: waveform_sig_loopback =5136;
21099: waveform_sig_loopback =4792;
21100: waveform_sig_loopback =3091;
21101: waveform_sig_loopback =5417;
21102: waveform_sig_loopback =4379;
21103: waveform_sig_loopback =3613;
21104: waveform_sig_loopback =4463;
21105: waveform_sig_loopback =4934;
21106: waveform_sig_loopback =3531;
21107: waveform_sig_loopback =3619;
21108: waveform_sig_loopback =5186;
21109: waveform_sig_loopback =4081;
21110: waveform_sig_loopback =2578;
21111: waveform_sig_loopback =4933;
21112: waveform_sig_loopback =4960;
21113: waveform_sig_loopback =2383;
21114: waveform_sig_loopback =3791;
21115: waveform_sig_loopback =5493;
21116: waveform_sig_loopback =2427;
21117: waveform_sig_loopback =5100;
21118: waveform_sig_loopback =3492;
21119: waveform_sig_loopback =510;
21120: waveform_sig_loopback =6600;
21121: waveform_sig_loopback =4026;
21122: waveform_sig_loopback =2700;
21123: waveform_sig_loopback =2609;
21124: waveform_sig_loopback =3316;
21125: waveform_sig_loopback =5336;
21126: waveform_sig_loopback =3073;
21127: waveform_sig_loopback =1864;
21128: waveform_sig_loopback =4494;
21129: waveform_sig_loopback =2705;
21130: waveform_sig_loopback =3858;
21131: waveform_sig_loopback =2796;
21132: waveform_sig_loopback =2486;
21133: waveform_sig_loopback =4639;
21134: waveform_sig_loopback =2015;
21135: waveform_sig_loopback =3068;
21136: waveform_sig_loopback =3308;
21137: waveform_sig_loopback =2902;
21138: waveform_sig_loopback =2310;
21139: waveform_sig_loopback =3621;
21140: waveform_sig_loopback =2848;
21141: waveform_sig_loopback =1797;
21142: waveform_sig_loopback =3621;
21143: waveform_sig_loopback =2640;
21144: waveform_sig_loopback =2219;
21145: waveform_sig_loopback =2499;
21146: waveform_sig_loopback =3489;
21147: waveform_sig_loopback =1790;
21148: waveform_sig_loopback =1833;
21149: waveform_sig_loopback =3821;
21150: waveform_sig_loopback =2080;
21151: waveform_sig_loopback =987;
21152: waveform_sig_loopback =3388;
21153: waveform_sig_loopback =3031;
21154: waveform_sig_loopback =748;
21155: waveform_sig_loopback =2132;
21156: waveform_sig_loopback =3684;
21157: waveform_sig_loopback =678;
21158: waveform_sig_loopback =3550;
21159: waveform_sig_loopback =1295;
21160: waveform_sig_loopback =-864;
21161: waveform_sig_loopback =4880;
21162: waveform_sig_loopback =1966;
21163: waveform_sig_loopback =1180;
21164: waveform_sig_loopback =644;
21165: waveform_sig_loopback =1797;
21166: waveform_sig_loopback =3650;
21167: waveform_sig_loopback =878;
21168: waveform_sig_loopback =514;
21169: waveform_sig_loopback =2531;
21170: waveform_sig_loopback =804;
21171: waveform_sig_loopback =2331;
21172: waveform_sig_loopback =566;
21173: waveform_sig_loopback =1028;
21174: waveform_sig_loopback =2719;
21175: waveform_sig_loopback =-65;
21176: waveform_sig_loopback =1607;
21177: waveform_sig_loopback =1168;
21178: waveform_sig_loopback =1132;
21179: waveform_sig_loopback =564;
21180: waveform_sig_loopback =1660;
21181: waveform_sig_loopback =1027;
21182: waveform_sig_loopback =-18;
21183: waveform_sig_loopback =1739;
21184: waveform_sig_loopback =796;
21185: waveform_sig_loopback =350;
21186: waveform_sig_loopback =658;
21187: waveform_sig_loopback =1708;
21188: waveform_sig_loopback =-150;
21189: waveform_sig_loopback =-36;
21190: waveform_sig_loopback =2171;
21191: waveform_sig_loopback =-115;
21192: waveform_sig_loopback =-749;
21193: waveform_sig_loopback =1750;
21194: waveform_sig_loopback =762;
21195: waveform_sig_loopback =-878;
21196: waveform_sig_loopback =249;
21197: waveform_sig_loopback =1646;
21198: waveform_sig_loopback =-950;
21199: waveform_sig_loopback =1491;
21200: waveform_sig_loopback =-693;
21201: waveform_sig_loopback =-2450;
21202: waveform_sig_loopback =2796;
21203: waveform_sig_loopback =256;
21204: waveform_sig_loopback =-875;
21205: waveform_sig_loopback =-1362;
21206: waveform_sig_loopback =283;
21207: waveform_sig_loopback =1431;
21208: waveform_sig_loopback =-1017;
21209: waveform_sig_loopback =-1164;
21210: waveform_sig_loopback =319;
21211: waveform_sig_loopback =-771;
21212: waveform_sig_loopback =312;
21213: waveform_sig_loopback =-1485;
21214: waveform_sig_loopback =-443;
21215: waveform_sig_loopback =439;
21216: waveform_sig_loopback =-1717;
21217: waveform_sig_loopback =-212;
21218: waveform_sig_loopback =-862;
21219: waveform_sig_loopback =-569;
21220: waveform_sig_loopback =-1450;
21221: waveform_sig_loopback =-117;
21222: waveform_sig_loopback =-933;
21223: waveform_sig_loopback =-1846;
21224: waveform_sig_loopback =-205;
21225: waveform_sig_loopback =-960;
21226: waveform_sig_loopback =-1670;
21227: waveform_sig_loopback =-1231;
21228: waveform_sig_loopback =28;
21229: waveform_sig_loopback =-2498;
21230: waveform_sig_loopback =-1550;
21231: waveform_sig_loopback =265;
21232: waveform_sig_loopback =-2376;
21233: waveform_sig_loopback =-2113;
21234: waveform_sig_loopback =-479;
21235: waveform_sig_loopback =-1109;
21236: waveform_sig_loopback =-2526;
21237: waveform_sig_loopback =-1988;
21238: waveform_sig_loopback =154;
21239: waveform_sig_loopback =-3091;
21240: waveform_sig_loopback =-377;
21241: waveform_sig_loopback =-2418;
21242: waveform_sig_loopback =-4593;
21243: waveform_sig_loopback =1235;
21244: waveform_sig_loopback =-1685;
21245: waveform_sig_loopback =-3118;
21246: waveform_sig_loopback =-2777;
21247: waveform_sig_loopback =-1690;
21248: waveform_sig_loopback =-544;
21249: waveform_sig_loopback =-2763;
21250: waveform_sig_loopback =-3220;
21251: waveform_sig_loopback =-1318;
21252: waveform_sig_loopback =-2657;
21253: waveform_sig_loopback =-1728;
21254: waveform_sig_loopback =-3145;
21255: waveform_sig_loopback =-2254;
21256: waveform_sig_loopback =-1584;
21257: waveform_sig_loopback =-3495;
21258: waveform_sig_loopback =-2051;
21259: waveform_sig_loopback =-2725;
21260: waveform_sig_loopback =-2415;
21261: waveform_sig_loopback =-3316;
21262: waveform_sig_loopback =-2018;
21263: waveform_sig_loopback =-2591;
21264: waveform_sig_loopback =-3890;
21265: waveform_sig_loopback =-1956;
21266: waveform_sig_loopback =-2634;
21267: waveform_sig_loopback =-3931;
21268: waveform_sig_loopback =-2393;
21269: waveform_sig_loopback =-2240;
21270: waveform_sig_loopback =-4326;
21271: waveform_sig_loopback =-2803;
21272: waveform_sig_loopback =-2226;
21273: waveform_sig_loopback =-3733;
21274: waveform_sig_loopback =-4062;
21275: waveform_sig_loopback =-2372;
21276: waveform_sig_loopback =-2504;
21277: waveform_sig_loopback =-4910;
21278: waveform_sig_loopback =-3236;
21279: waveform_sig_loopback =-1722;
21280: waveform_sig_loopback =-5185;
21281: waveform_sig_loopback =-1606;
21282: waveform_sig_loopback =-4793;
21283: waveform_sig_loopback =-5963;
21284: waveform_sig_loopback =-376;
21285: waveform_sig_loopback =-3793;
21286: waveform_sig_loopback =-4617;
21287: waveform_sig_loopback =-4582;
21288: waveform_sig_loopback =-3344;
21289: waveform_sig_loopback =-2259;
21290: waveform_sig_loopback =-4506;
21291: waveform_sig_loopback =-4880;
21292: waveform_sig_loopback =-3038;
21293: waveform_sig_loopback =-4266;
21294: waveform_sig_loopback =-3583;
21295: waveform_sig_loopback =-4707;
21296: waveform_sig_loopback =-3950;
21297: waveform_sig_loopback =-3408;
21298: waveform_sig_loopback =-4878;
21299: waveform_sig_loopback =-4056;
21300: waveform_sig_loopback =-4212;
21301: waveform_sig_loopback =-3878;
21302: waveform_sig_loopback =-5429;
21303: waveform_sig_loopback =-3042;
21304: waveform_sig_loopback =-4672;
21305: waveform_sig_loopback =-5380;
21306: waveform_sig_loopback =-3109;
21307: waveform_sig_loopback =-4950;
21308: waveform_sig_loopback =-5039;
21309: waveform_sig_loopback =-4115;
21310: waveform_sig_loopback =-4000;
21311: waveform_sig_loopback =-5508;
21312: waveform_sig_loopback =-4820;
21313: waveform_sig_loopback =-3518;
21314: waveform_sig_loopback =-5249;
21315: waveform_sig_loopback =-5864;
21316: waveform_sig_loopback =-3542;
21317: waveform_sig_loopback =-4304;
21318: waveform_sig_loopback =-6460;
21319: waveform_sig_loopback =-4504;
21320: waveform_sig_loopback =-3446;
21321: waveform_sig_loopback =-6600;
21322: waveform_sig_loopback =-2973;
21323: waveform_sig_loopback =-6572;
21324: waveform_sig_loopback =-7209;
21325: waveform_sig_loopback =-1772;
21326: waveform_sig_loopback =-5455;
21327: waveform_sig_loopback =-6061;
21328: waveform_sig_loopback =-5962;
21329: waveform_sig_loopback =-4923;
21330: waveform_sig_loopback =-3490;
21331: waveform_sig_loopback =-6184;
21332: waveform_sig_loopback =-6367;
21333: waveform_sig_loopback =-4147;
21334: waveform_sig_loopback =-5999;
21335: waveform_sig_loopback =-4775;
21336: waveform_sig_loopback =-6112;
21337: waveform_sig_loopback =-5599;
21338: waveform_sig_loopback =-4397;
21339: waveform_sig_loopback =-6445;
21340: waveform_sig_loopback =-5467;
21341: waveform_sig_loopback =-5201;
21342: waveform_sig_loopback =-5723;
21343: waveform_sig_loopback =-6395;
21344: waveform_sig_loopback =-4337;
21345: waveform_sig_loopback =-6471;
21346: waveform_sig_loopback =-6156;
21347: waveform_sig_loopback =-4894;
21348: waveform_sig_loopback =-6104;
21349: waveform_sig_loopback =-6149;
21350: waveform_sig_loopback =-5794;
21351: waveform_sig_loopback =-4976;
21352: waveform_sig_loopback =-7012;
21353: waveform_sig_loopback =-5976;
21354: waveform_sig_loopback =-4670;
21355: waveform_sig_loopback =-6799;
21356: waveform_sig_loopback =-6856;
21357: waveform_sig_loopback =-4850;
21358: waveform_sig_loopback =-5592;
21359: waveform_sig_loopback =-7759;
21360: waveform_sig_loopback =-5521;
21361: waveform_sig_loopback =-4815;
21362: waveform_sig_loopback =-8064;
21363: waveform_sig_loopback =-3749;
21364: waveform_sig_loopback =-8252;
21365: waveform_sig_loopback =-7918;
21366: waveform_sig_loopback =-3154;
21367: waveform_sig_loopback =-7000;
21368: waveform_sig_loopback =-6562;
21369: waveform_sig_loopback =-7506;
21370: waveform_sig_loopback =-5964;
21371: waveform_sig_loopback =-4466;
21372: waveform_sig_loopback =-7654;
21373: waveform_sig_loopback =-6904;
21374: waveform_sig_loopback =-5590;
21375: waveform_sig_loopback =-7181;
21376: waveform_sig_loopback =-5337;
21377: waveform_sig_loopback =-7705;
21378: waveform_sig_loopback =-6295;
21379: waveform_sig_loopback =-5500;
21380: waveform_sig_loopback =-7784;
21381: waveform_sig_loopback =-5985;
21382: waveform_sig_loopback =-6720;
21383: waveform_sig_loopback =-6620;
21384: waveform_sig_loopback =-7108;
21385: waveform_sig_loopback =-5686;
21386: waveform_sig_loopback =-7222;
21387: waveform_sig_loopback =-7168;
21388: waveform_sig_loopback =-5789;
21389: waveform_sig_loopback =-7005;
21390: waveform_sig_loopback =-7203;
21391: waveform_sig_loopback =-6502;
21392: waveform_sig_loopback =-5947;
21393: waveform_sig_loopback =-7946;
21394: waveform_sig_loopback =-6888;
21395: waveform_sig_loopback =-5339;
21396: waveform_sig_loopback =-7910;
21397: waveform_sig_loopback =-7666;
21398: waveform_sig_loopback =-5371;
21399: waveform_sig_loopback =-6813;
21400: waveform_sig_loopback =-8257;
21401: waveform_sig_loopback =-6302;
21402: waveform_sig_loopback =-5922;
21403: waveform_sig_loopback =-8164;
21404: waveform_sig_loopback =-4920;
21405: waveform_sig_loopback =-9149;
21406: waveform_sig_loopback =-8194;
21407: waveform_sig_loopback =-4156;
21408: waveform_sig_loopback =-7330;
21409: waveform_sig_loopback =-7720;
21410: waveform_sig_loopback =-8275;
21411: waveform_sig_loopback =-5995;
21412: waveform_sig_loopback =-5611;
21413: waveform_sig_loopback =-8342;
21414: waveform_sig_loopback =-7383;
21415: waveform_sig_loopback =-6493;
21416: waveform_sig_loopback =-7428;
21417: waveform_sig_loopback =-6285;
21418: waveform_sig_loopback =-8425;
21419: waveform_sig_loopback =-6387;
21420: waveform_sig_loopback =-6574;
21421: waveform_sig_loopback =-8193;
21422: waveform_sig_loopback =-6473;
21423: waveform_sig_loopback =-7413;
21424: waveform_sig_loopback =-6954;
21425: waveform_sig_loopback =-7827;
21426: waveform_sig_loopback =-6144;
21427: waveform_sig_loopback =-7695;
21428: waveform_sig_loopback =-7717;
21429: waveform_sig_loopback =-6342;
21430: waveform_sig_loopback =-7293;
21431: waveform_sig_loopback =-7843;
21432: waveform_sig_loopback =-6884;
21433: waveform_sig_loopback =-6325;
21434: waveform_sig_loopback =-8591;
21435: waveform_sig_loopback =-6957;
21436: waveform_sig_loopback =-5955;
21437: waveform_sig_loopback =-8371;
21438: waveform_sig_loopback =-7689;
21439: waveform_sig_loopback =-5995;
21440: waveform_sig_loopback =-7156;
21441: waveform_sig_loopback =-8479;
21442: waveform_sig_loopback =-6727;
21443: waveform_sig_loopback =-6075;
21444: waveform_sig_loopback =-8474;
21445: waveform_sig_loopback =-5405;
21446: waveform_sig_loopback =-9250;
21447: waveform_sig_loopback =-8519;
21448: waveform_sig_loopback =-4336;
21449: waveform_sig_loopback =-7465;
21450: waveform_sig_loopback =-8316;
21451: waveform_sig_loopback =-8044;
21452: waveform_sig_loopback =-6364;
21453: waveform_sig_loopback =-5937;
21454: waveform_sig_loopback =-8203;
21455: waveform_sig_loopback =-7843;
21456: waveform_sig_loopback =-6468;
21457: waveform_sig_loopback =-7518;
21458: waveform_sig_loopback =-6685;
21459: waveform_sig_loopback =-8273;
21460: waveform_sig_loopback =-6586;
21461: waveform_sig_loopback =-6753;
21462: waveform_sig_loopback =-8086;
21463: waveform_sig_loopback =-6684;
21464: waveform_sig_loopback =-7336;
21465: waveform_sig_loopback =-7036;
21466: waveform_sig_loopback =-7827;
21467: waveform_sig_loopback =-6103;
21468: waveform_sig_loopback =-7679;
21469: waveform_sig_loopback =-7801;
21470: waveform_sig_loopback =-6159;
21471: waveform_sig_loopback =-7297;
21472: waveform_sig_loopback =-8013;
21473: waveform_sig_loopback =-6394;
21474: waveform_sig_loopback =-6671;
21475: waveform_sig_loopback =-8416;
21476: waveform_sig_loopback =-6601;
21477: waveform_sig_loopback =-6216;
21478: waveform_sig_loopback =-8003;
21479: waveform_sig_loopback =-7657;
21480: waveform_sig_loopback =-5841;
21481: waveform_sig_loopback =-6882;
21482: waveform_sig_loopback =-8590;
21483: waveform_sig_loopback =-6313;
21484: waveform_sig_loopback =-5933;
21485: waveform_sig_loopback =-8452;
21486: waveform_sig_loopback =-4922;
21487: waveform_sig_loopback =-9366;
21488: waveform_sig_loopback =-8123;
21489: waveform_sig_loopback =-3908;
21490: waveform_sig_loopback =-7509;
21491: waveform_sig_loopback =-8035;
21492: waveform_sig_loopback =-7578;
21493: waveform_sig_loopback =-6262;
21494: waveform_sig_loopback =-5470;
21495: waveform_sig_loopback =-8043;
21496: waveform_sig_loopback =-7580;
21497: waveform_sig_loopback =-5902;
21498: waveform_sig_loopback =-7376;
21499: waveform_sig_loopback =-6244;
21500: waveform_sig_loopback =-7798;
21501: waveform_sig_loopback =-6331;
21502: waveform_sig_loopback =-6273;
21503: waveform_sig_loopback =-7658;
21504: waveform_sig_loopback =-6372;
21505: waveform_sig_loopback =-6752;
21506: waveform_sig_loopback =-6700;
21507: waveform_sig_loopback =-7392;
21508: waveform_sig_loopback =-5460;
21509: waveform_sig_loopback =-7448;
21510: waveform_sig_loopback =-7192;
21511: waveform_sig_loopback =-5557;
21512: waveform_sig_loopback =-7036;
21513: waveform_sig_loopback =-7301;
21514: waveform_sig_loopback =-5810;
21515: waveform_sig_loopback =-6323;
21516: waveform_sig_loopback =-7635;
21517: waveform_sig_loopback =-6162;
21518: waveform_sig_loopback =-5685;
21519: waveform_sig_loopback =-7285;
21520: waveform_sig_loopback =-7256;
21521: waveform_sig_loopback =-5076;
21522: waveform_sig_loopback =-6316;
21523: waveform_sig_loopback =-8144;
21524: waveform_sig_loopback =-5272;
21525: waveform_sig_loopback =-5593;
21526: waveform_sig_loopback =-7762;
21527: waveform_sig_loopback =-3969;
21528: waveform_sig_loopback =-9199;
21529: waveform_sig_loopback =-6897;
21530: waveform_sig_loopback =-3265;
21531: waveform_sig_loopback =-7126;
21532: waveform_sig_loopback =-6921;
21533: waveform_sig_loopback =-7020;
21534: waveform_sig_loopback =-5431;
21535: waveform_sig_loopback =-4572;
21536: waveform_sig_loopback =-7598;
21537: waveform_sig_loopback =-6444;
21538: waveform_sig_loopback =-5186;
21539: waveform_sig_loopback =-6667;
21540: waveform_sig_loopback =-5240;
21541: waveform_sig_loopback =-7162;
21542: waveform_sig_loopback =-5353;
21543: waveform_sig_loopback =-5396;
21544: waveform_sig_loopback =-6885;
21545: waveform_sig_loopback =-5464;
21546: waveform_sig_loopback =-5789;
21547: waveform_sig_loopback =-5927;
21548: waveform_sig_loopback =-6436;
21549: waveform_sig_loopback =-4423;
21550: waveform_sig_loopback =-6777;
21551: waveform_sig_loopback =-5937;
21552: waveform_sig_loopback =-4683;
21553: waveform_sig_loopback =-6288;
21554: waveform_sig_loopback =-5905;
21555: waveform_sig_loopback =-5108;
21556: waveform_sig_loopback =-5289;
21557: waveform_sig_loopback =-6476;
21558: waveform_sig_loopback =-5397;
21559: waveform_sig_loopback =-4270;
21560: waveform_sig_loopback =-6623;
21561: waveform_sig_loopback =-6088;
21562: waveform_sig_loopback =-3670;
21563: waveform_sig_loopback =-5775;
21564: waveform_sig_loopback =-6750;
21565: waveform_sig_loopback =-4117;
21566: waveform_sig_loopback =-4833;
21567: waveform_sig_loopback =-6262;
21568: waveform_sig_loopback =-3066;
21569: waveform_sig_loopback =-8221;
21570: waveform_sig_loopback =-5347;
21571: waveform_sig_loopback =-2408;
21572: waveform_sig_loopback =-5900;
21573: waveform_sig_loopback =-5725;
21574: waveform_sig_loopback =-6035;
21575: waveform_sig_loopback =-3933;
21576: waveform_sig_loopback =-3446;
21577: waveform_sig_loopback =-6656;
21578: waveform_sig_loopback =-4854;
21579: waveform_sig_loopback =-4216;
21580: waveform_sig_loopback =-5345;
21581: waveform_sig_loopback =-3888;
21582: waveform_sig_loopback =-6154;
21583: waveform_sig_loopback =-3784;
21584: waveform_sig_loopback =-4274;
21585: waveform_sig_loopback =-5663;
21586: waveform_sig_loopback =-3996;
21587: waveform_sig_loopback =-4585;
21588: waveform_sig_loopback =-4755;
21589: waveform_sig_loopback =-4806;
21590: waveform_sig_loopback =-3325;
21591: waveform_sig_loopback =-5528;
21592: waveform_sig_loopback =-4264;
21593: waveform_sig_loopback =-3727;
21594: waveform_sig_loopback =-4668;
21595: waveform_sig_loopback =-4666;
21596: waveform_sig_loopback =-3854;
21597: waveform_sig_loopback =-3590;
21598: waveform_sig_loopback =-5495;
21599: waveform_sig_loopback =-3669;
21600: waveform_sig_loopback =-2885;
21601: waveform_sig_loopback =-5496;
21602: waveform_sig_loopback =-4267;
21603: waveform_sig_loopback =-2461;
21604: waveform_sig_loopback =-4399;
21605: waveform_sig_loopback =-5081;
21606: waveform_sig_loopback =-2779;
21607: waveform_sig_loopback =-3364;
21608: waveform_sig_loopback =-4640;
21609: waveform_sig_loopback =-1794;
21610: waveform_sig_loopback =-6758;
21611: waveform_sig_loopback =-3593;
21612: waveform_sig_loopback =-1042;
21613: waveform_sig_loopback =-4375;
21614: waveform_sig_loopback =-4248;
21615: waveform_sig_loopback =-4487;
21616: waveform_sig_loopback =-2182;
21617: waveform_sig_loopback =-2163;
21618: waveform_sig_loopback =-5123;
21619: waveform_sig_loopback =-3010;
21620: waveform_sig_loopback =-3021;
21621: waveform_sig_loopback =-3483;
21622: waveform_sig_loopback =-2386;
21623: waveform_sig_loopback =-4771;
21624: waveform_sig_loopback =-1755;
21625: waveform_sig_loopback =-3088;
21626: waveform_sig_loopback =-3917;
21627: waveform_sig_loopback =-2230;
21628: waveform_sig_loopback =-3261;
21629: waveform_sig_loopback =-2844;
21630: waveform_sig_loopback =-3226;
21631: waveform_sig_loopback =-1882;
21632: waveform_sig_loopback =-3560;
21633: waveform_sig_loopback =-2896;
21634: waveform_sig_loopback =-1964;
21635: waveform_sig_loopback =-2899;
21636: waveform_sig_loopback =-3314;
21637: waveform_sig_loopback =-1771;
21638: waveform_sig_loopback =-2170;
21639: waveform_sig_loopback =-3821;
21640: waveform_sig_loopback =-1716;
21641: waveform_sig_loopback =-1467;
21642: waveform_sig_loopback =-3712;
21643: waveform_sig_loopback =-2454;
21644: waveform_sig_loopback =-818;
21645: waveform_sig_loopback =-2748;
21646: waveform_sig_loopback =-3304;
21647: waveform_sig_loopback =-1078;
21648: waveform_sig_loopback =-1705;
21649: waveform_sig_loopback =-2734;
21650: waveform_sig_loopback =-291;
21651: waveform_sig_loopback =-4906;
21652: waveform_sig_loopback =-1727;
21653: waveform_sig_loopback =510;
21654: waveform_sig_loopback =-2282;
21655: waveform_sig_loopback =-2920;
21656: waveform_sig_loopback =-2473;
21657: waveform_sig_loopback =-247;
21658: waveform_sig_loopback =-707;
21659: waveform_sig_loopback =-3036;
21660: waveform_sig_loopback =-1422;
21661: waveform_sig_loopback =-1195;
21662: waveform_sig_loopback =-1363;
21663: waveform_sig_loopback =-1080;
21664: waveform_sig_loopback =-2563;
21665: waveform_sig_loopback =16;
21666: waveform_sig_loopback =-1559;
21667: waveform_sig_loopback =-1672;
21668: waveform_sig_loopback =-771;
21669: waveform_sig_loopback =-1249;
21670: waveform_sig_loopback =-1055;
21671: waveform_sig_loopback =-1530;
21672: waveform_sig_loopback =185;
21673: waveform_sig_loopback =-1954;
21674: waveform_sig_loopback =-953;
21675: waveform_sig_loopback =-109;
21676: waveform_sig_loopback =-1125;
21677: waveform_sig_loopback =-1491;
21678: waveform_sig_loopback =178;
21679: waveform_sig_loopback =-432;
21680: waveform_sig_loopback =-2027;
21681: waveform_sig_loopback =408;
21682: waveform_sig_loopback =83;
21683: waveform_sig_loopback =-1745;
21684: waveform_sig_loopback =-415;
21685: waveform_sig_loopback =726;
21686: waveform_sig_loopback =-604;
21687: waveform_sig_loopback =-1619;
21688: waveform_sig_loopback =921;
21689: waveform_sig_loopback =252;
21690: waveform_sig_loopback =-1080;
21691: waveform_sig_loopback =1838;
21692: waveform_sig_loopback =-3212;
21693: waveform_sig_loopback =268;
21694: waveform_sig_loopback =2597;
21695: waveform_sig_loopback =-814;
21696: waveform_sig_loopback =-916;
21697: waveform_sig_loopback =-279;
21698: waveform_sig_loopback =1277;
21699: waveform_sig_loopback =1321;
21700: waveform_sig_loopback =-1191;
21701: waveform_sig_loopback =362;
21702: waveform_sig_loopback =936;
21703: waveform_sig_loopback =236;
21704: waveform_sig_loopback =894;
21705: waveform_sig_loopback =-513;
21706: waveform_sig_loopback =1599;
21707: waveform_sig_loopback =467;
21708: waveform_sig_loopback =215;
21709: waveform_sig_loopback =1063;
21710: waveform_sig_loopback =728;
21711: waveform_sig_loopback =496;
21712: waveform_sig_loopback =554;
21713: waveform_sig_loopback =2215;
21714: waveform_sig_loopback =-264;
21715: waveform_sig_loopback =748;
21716: waveform_sig_loopback =2020;
21717: waveform_sig_loopback =748;
21718: waveform_sig_loopback =495;
21719: waveform_sig_loopback =2084;
21720: waveform_sig_loopback =1072;
21721: waveform_sig_loopback =410;
21722: waveform_sig_loopback =2159;
21723: waveform_sig_loopback =1679;
21724: waveform_sig_loopback =442;
21725: waveform_sig_loopback =1301;
21726: waveform_sig_loopback =2792;
21727: waveform_sig_loopback =1174;
21728: waveform_sig_loopback =45;
21729: waveform_sig_loopback =3398;
21730: waveform_sig_loopback =1624;
21731: waveform_sig_loopback =819;
21732: waveform_sig_loopback =4008;
21733: waveform_sig_loopback =-1873;
21734: waveform_sig_loopback =2725;
21735: waveform_sig_loopback =4163;
21736: waveform_sig_loopback =862;
21737: waveform_sig_loopback =1319;
21738: waveform_sig_loopback =1303;
21739: waveform_sig_loopback =3274;
21740: waveform_sig_loopback =3103;
21741: waveform_sig_loopback =516;
21742: waveform_sig_loopback =2451;
21743: waveform_sig_loopback =2624;
21744: waveform_sig_loopback =2071;
21745: waveform_sig_loopback =2741;
21746: waveform_sig_loopback =1366;
21747: waveform_sig_loopback =3377;
21748: waveform_sig_loopback =2337;
21749: waveform_sig_loopback =2120;
21750: waveform_sig_loopback =2697;
21751: waveform_sig_loopback =2855;
21752: waveform_sig_loopback =2329;
21753: waveform_sig_loopback =2230;
21754: waveform_sig_loopback =4168;
21755: waveform_sig_loopback =1194;
21756: waveform_sig_loopback =3311;
21757: waveform_sig_loopback =3491;
21758: waveform_sig_loopback =2100;
21759: waveform_sig_loopback =2916;
21760: waveform_sig_loopback =3499;
21761: waveform_sig_loopback =3076;
21762: waveform_sig_loopback =2069;
21763: waveform_sig_loopback =3833;
21764: waveform_sig_loopback =3870;
21765: waveform_sig_loopback =1765;
21766: waveform_sig_loopback =3268;
21767: waveform_sig_loopback =4626;
21768: waveform_sig_loopback =2671;
21769: waveform_sig_loopback =2066;
21770: waveform_sig_loopback =5043;
21771: waveform_sig_loopback =3257;
21772: waveform_sig_loopback =2889;
21773: waveform_sig_loopback =5467;
21774: waveform_sig_loopback =-243;
21775: waveform_sig_loopback =4805;
21776: waveform_sig_loopback =5758;
21777: waveform_sig_loopback =2471;
21778: waveform_sig_loopback =3092;
21779: waveform_sig_loopback =3002;
21780: waveform_sig_loopback =5131;
21781: waveform_sig_loopback =4815;
21782: waveform_sig_loopback =1983;
21783: waveform_sig_loopback =4451;
21784: waveform_sig_loopback =4233;
21785: waveform_sig_loopback =3710;
21786: waveform_sig_loopback =4589;
21787: waveform_sig_loopback =2824;
21788: waveform_sig_loopback =5231;
21789: waveform_sig_loopback =4066;
21790: waveform_sig_loopback =3493;
21791: waveform_sig_loopback =4620;
21792: waveform_sig_loopback =4418;
21793: waveform_sig_loopback =3686;
21794: waveform_sig_loopback =4417;
21795: waveform_sig_loopback =5293;
21796: waveform_sig_loopback =2975;
21797: waveform_sig_loopback =5115;
21798: waveform_sig_loopback =4710;
21799: waveform_sig_loopback =4161;
21800: waveform_sig_loopback =4171;
21801: waveform_sig_loopback =5240;
21802: waveform_sig_loopback =4777;
21803: waveform_sig_loopback =3314;
21804: waveform_sig_loopback =5703;
21805: waveform_sig_loopback =5261;
21806: waveform_sig_loopback =3299;
21807: waveform_sig_loopback =4980;
21808: waveform_sig_loopback =6175;
21809: waveform_sig_loopback =4089;
21810: waveform_sig_loopback =3698;
21811: waveform_sig_loopback =6731;
21812: waveform_sig_loopback =4401;
21813: waveform_sig_loopback =4864;
21814: waveform_sig_loopback =6686;
21815: waveform_sig_loopback =1152;
21816: waveform_sig_loopback =6850;
21817: waveform_sig_loopback =6718;
21818: waveform_sig_loopback =4178;
21819: waveform_sig_loopback =4594;
21820: waveform_sig_loopback =4294;
21821: waveform_sig_loopback =7024;
21822: waveform_sig_loopback =5853;
21823: waveform_sig_loopback =3446;
21824: waveform_sig_loopback =6222;
21825: waveform_sig_loopback =5158;
21826: waveform_sig_loopback =5489;
21827: waveform_sig_loopback =5854;
21828: waveform_sig_loopback =4062;
21829: waveform_sig_loopback =7066;
21830: waveform_sig_loopback =4964;
21831: waveform_sig_loopback =5035;
21832: waveform_sig_loopback =6196;
21833: waveform_sig_loopback =5385;
21834: waveform_sig_loopback =5348;
21835: waveform_sig_loopback =5706;
21836: waveform_sig_loopback =6459;
21837: waveform_sig_loopback =4583;
21838: waveform_sig_loopback =6185;
21839: waveform_sig_loopback =6144;
21840: waveform_sig_loopback =5404;
21841: waveform_sig_loopback =5408;
21842: waveform_sig_loopback =6664;
21843: waveform_sig_loopback =5852;
21844: waveform_sig_loopback =4677;
21845: waveform_sig_loopback =7025;
21846: waveform_sig_loopback =6445;
21847: waveform_sig_loopback =4411;
21848: waveform_sig_loopback =6440;
21849: waveform_sig_loopback =7329;
21850: waveform_sig_loopback =5062;
21851: waveform_sig_loopback =5272;
21852: waveform_sig_loopback =7640;
21853: waveform_sig_loopback =5601;
21854: waveform_sig_loopback =6329;
21855: waveform_sig_loopback =7283;
21856: waveform_sig_loopback =2743;
21857: waveform_sig_loopback =7902;
21858: waveform_sig_loopback =7626;
21859: waveform_sig_loopback =5689;
21860: waveform_sig_loopback =5131;
21861: waveform_sig_loopback =5815;
21862: waveform_sig_loopback =8123;
21863: waveform_sig_loopback =6511;
21864: waveform_sig_loopback =5034;
21865: waveform_sig_loopback =6933;
21866: waveform_sig_loopback =6274;
21867: waveform_sig_loopback =6838;
21868: waveform_sig_loopback =6386;
21869: waveform_sig_loopback =5470;
21870: waveform_sig_loopback =7999;
21871: waveform_sig_loopback =5778;
21872: waveform_sig_loopback =6378;
21873: waveform_sig_loopback =6843;
21874: waveform_sig_loopback =6536;
21875: waveform_sig_loopback =6304;
21876: waveform_sig_loopback =6621;
21877: waveform_sig_loopback =7412;
21878: waveform_sig_loopback =5520;
21879: waveform_sig_loopback =7089;
21880: waveform_sig_loopback =7080;
21881: waveform_sig_loopback =6423;
21882: waveform_sig_loopback =6091;
21883: waveform_sig_loopback =7870;
21884: waveform_sig_loopback =6530;
21885: waveform_sig_loopback =5519;
21886: waveform_sig_loopback =8258;
21887: waveform_sig_loopback =6820;
21888: waveform_sig_loopback =5517;
21889: waveform_sig_loopback =7358;
21890: waveform_sig_loopback =7876;
21891: waveform_sig_loopback =6080;
21892: waveform_sig_loopback =5945;
21893: waveform_sig_loopback =8422;
21894: waveform_sig_loopback =6544;
21895: waveform_sig_loopback =6850;
21896: waveform_sig_loopback =8070;
21897: waveform_sig_loopback =3606;
21898: waveform_sig_loopback =8481;
21899: waveform_sig_loopback =8664;
21900: waveform_sig_loopback =6064;
21901: waveform_sig_loopback =5843;
21902: waveform_sig_loopback =6871;
21903: waveform_sig_loopback =8375;
21904: waveform_sig_loopback =7424;
21905: waveform_sig_loopback =5609;
21906: waveform_sig_loopback =7485;
21907: waveform_sig_loopback =7088;
21908: waveform_sig_loopback =7290;
21909: waveform_sig_loopback =6952;
21910: waveform_sig_loopback =6275;
21911: waveform_sig_loopback =8391;
21912: waveform_sig_loopback =6352;
21913: waveform_sig_loopback =7066;
21914: waveform_sig_loopback =7233;
21915: waveform_sig_loopback =7192;
21916: waveform_sig_loopback =6805;
21917: waveform_sig_loopback =7096;
21918: waveform_sig_loopback =8059;
21919: waveform_sig_loopback =5897;
21920: waveform_sig_loopback =7547;
21921: waveform_sig_loopback =7769;
21922: waveform_sig_loopback =6533;
21923: waveform_sig_loopback =6726;
21924: waveform_sig_loopback =8409;
21925: waveform_sig_loopback =6547;
21926: waveform_sig_loopback =6283;
21927: waveform_sig_loopback =8496;
21928: waveform_sig_loopback =7071;
21929: waveform_sig_loopback =6103;
21930: waveform_sig_loopback =7543;
21931: waveform_sig_loopback =8264;
21932: waveform_sig_loopback =6484;
21933: waveform_sig_loopback =6031;
21934: waveform_sig_loopback =9086;
21935: waveform_sig_loopback =6525;
21936: waveform_sig_loopback =7201;
21937: waveform_sig_loopback =8518;
21938: waveform_sig_loopback =3456;
21939: waveform_sig_loopback =9178;
21940: waveform_sig_loopback =8788;
21941: waveform_sig_loopback =5949;
21942: waveform_sig_loopback =6431;
21943: waveform_sig_loopback =6943;
21944: waveform_sig_loopback =8566;
21945: waveform_sig_loopback =7716;
21946: waveform_sig_loopback =5578;
21947: waveform_sig_loopback =7851;
21948: waveform_sig_loopback =7267;
21949: waveform_sig_loopback =7257;
21950: waveform_sig_loopback =7233;
21951: waveform_sig_loopback =6409;
21952: waveform_sig_loopback =8364;
21953: waveform_sig_loopback =6626;
21954: waveform_sig_loopback =7023;
21955: waveform_sig_loopback =7280;
21956: waveform_sig_loopback =7457;
21957: waveform_sig_loopback =6609;
21958: waveform_sig_loopback =7308;
21959: waveform_sig_loopback =8015;
21960: waveform_sig_loopback =5663;
21961: waveform_sig_loopback =7948;
21962: waveform_sig_loopback =7641;
21963: waveform_sig_loopback =6263;
21964: waveform_sig_loopback =7097;
21965: waveform_sig_loopback =8057;
21966: waveform_sig_loopback =6610;
21967: waveform_sig_loopback =6423;
21968: waveform_sig_loopback =8011;
21969: waveform_sig_loopback =7300;
21970: waveform_sig_loopback =5841;
21971: waveform_sig_loopback =7443;
21972: waveform_sig_loopback =8350;
21973: waveform_sig_loopback =5919;
21974: waveform_sig_loopback =6194;
21975: waveform_sig_loopback =9023;
21976: waveform_sig_loopback =5976;
21977: waveform_sig_loopback =7497;
21978: waveform_sig_loopback =7972;
21979: waveform_sig_loopback =3182;
21980: waveform_sig_loopback =9442;
21981: waveform_sig_loopback =8136;
21982: waveform_sig_loopback =5781;
21983: waveform_sig_loopback =6259;
21984: waveform_sig_loopback =6407;
21985: waveform_sig_loopback =8606;
21986: waveform_sig_loopback =7216;
21987: waveform_sig_loopback =5065;
21988: waveform_sig_loopback =7893;
21989: waveform_sig_loopback =6659;
21990: waveform_sig_loopback =7055;
21991: waveform_sig_loopback =6897;
21992: waveform_sig_loopback =5873;
21993: waveform_sig_loopback =8241;
21994: waveform_sig_loopback =6108;
21995: waveform_sig_loopback =6586;
21996: waveform_sig_loopback =7055;
21997: waveform_sig_loopback =6936;
21998: waveform_sig_loopback =6063;
21999: waveform_sig_loopback =7109;
22000: waveform_sig_loopback =7440;
22001: waveform_sig_loopback =5249;
22002: waveform_sig_loopback =7648;
22003: waveform_sig_loopback =6782;
22004: waveform_sig_loopback =5961;
22005: waveform_sig_loopback =6633;
22006: waveform_sig_loopback =7350;
22007: waveform_sig_loopback =6201;
22008: waveform_sig_loopback =5714;
22009: waveform_sig_loopback =7520;
22010: waveform_sig_loopback =6888;
22011: waveform_sig_loopback =4879;
22012: waveform_sig_loopback =7165;
22013: waveform_sig_loopback =7710;
22014: waveform_sig_loopback =4951;
22015: waveform_sig_loopback =6098;
22016: waveform_sig_loopback =7986;
22017: waveform_sig_loopback =5347;
22018: waveform_sig_loopback =7168;
22019: waveform_sig_loopback =6726;
22020: waveform_sig_loopback =3003;
22021: waveform_sig_loopback =8637;
22022: waveform_sig_loopback =7299;
22023: waveform_sig_loopback =5365;
22024: waveform_sig_loopback =5241;
22025: waveform_sig_loopback =5896;
22026: waveform_sig_loopback =7920;
22027: waveform_sig_loopback =6276;
22028: waveform_sig_loopback =4396;
22029: waveform_sig_loopback =7128;
22030: waveform_sig_loopback =5704;
22031: waveform_sig_loopback =6459;
22032: waveform_sig_loopback =5935;
22033: waveform_sig_loopback =5000;
22034: waveform_sig_loopback =7590;
22035: waveform_sig_loopback =5053;
22036: waveform_sig_loopback =5783;
22037: waveform_sig_loopback =6307;
22038: waveform_sig_loopback =5797;
22039: waveform_sig_loopback =5301;
22040: waveform_sig_loopback =6378;
22041: waveform_sig_loopback =6082;
22042: waveform_sig_loopback =4685;
22043: waveform_sig_loopback =6484;
22044: waveform_sig_loopback =5789;
22045: waveform_sig_loopback =5305;
22046: waveform_sig_loopback =5299;
22047: waveform_sig_loopback =6653;
22048: waveform_sig_loopback =5084;
22049: waveform_sig_loopback =4577;
22050: waveform_sig_loopback =6970;
22051: waveform_sig_loopback =5422;
22052: waveform_sig_loopback =3985;
22053: waveform_sig_loopback =6375;
22054: waveform_sig_loopback =6262;
22055: waveform_sig_loopback =4186;
22056: waveform_sig_loopback =4904;
22057: waveform_sig_loopback =6903;
22058: waveform_sig_loopback =4232;
22059: waveform_sig_loopback =5939;
22060: waveform_sig_loopback =5643;
22061: waveform_sig_loopback =1948;
22062: waveform_sig_loopback =7491;
22063: waveform_sig_loopback =5868;
22064: waveform_sig_loopback =4382;
22065: waveform_sig_loopback =4066;
22066: waveform_sig_loopback =4754;
22067: waveform_sig_loopback =6670;
22068: waveform_sig_loopback =4966;
22069: waveform_sig_loopback =3515;
22070: waveform_sig_loopback =5747;
22071: waveform_sig_loopback =4302;
22072: waveform_sig_loopback =5567;
22073: waveform_sig_loopback =4409;
22074: waveform_sig_loopback =3887;
22075: waveform_sig_loopback =6352;
22076: waveform_sig_loopback =3486;
22077: waveform_sig_loopback =4884;
22078: waveform_sig_loopback =4750;
22079: waveform_sig_loopback =4382;
22080: waveform_sig_loopback =4345;
22081: waveform_sig_loopback =4706;
22082: waveform_sig_loopback =4869;
22083: waveform_sig_loopback =3398;
22084: waveform_sig_loopback =4914;
22085: waveform_sig_loopback =4784;
22086: waveform_sig_loopback =3506;
22087: waveform_sig_loopback =4077;
22088: waveform_sig_loopback =5485;
22089: waveform_sig_loopback =3260;
22090: waveform_sig_loopback =3507;
22091: waveform_sig_loopback =5476;
22092: waveform_sig_loopback =3879;
22093: waveform_sig_loopback =2767;
22094: waveform_sig_loopback =4797;
22095: waveform_sig_loopback =4853;
22096: waveform_sig_loopback =2728;
22097: waveform_sig_loopback =3474;
22098: waveform_sig_loopback =5436;
22099: waveform_sig_loopback =2798;
22100: waveform_sig_loopback =4692;
22101: waveform_sig_loopback =3675;
22102: waveform_sig_loopback =618;
22103: waveform_sig_loopback =6182;
22104: waveform_sig_loopback =4409;
22105: waveform_sig_loopback =2660;
22106: waveform_sig_loopback =2321;
22107: waveform_sig_loopback =3709;
22108: waveform_sig_loopback =5027;
22109: waveform_sig_loopback =3098;
22110: waveform_sig_loopback =2184;
22111: waveform_sig_loopback =4027;
22112: waveform_sig_loopback =3045;
22113: waveform_sig_loopback =3813;
22114: waveform_sig_loopback =2504;
22115: waveform_sig_loopback =2931;
22116: waveform_sig_loopback =4268;
22117: waveform_sig_loopback =1982;
22118: waveform_sig_loopback =3416;
22119: waveform_sig_loopback =2807;
22120: waveform_sig_loopback =3259;
22121: waveform_sig_loopback =2211;
22122: waveform_sig_loopback =3266;
22123: waveform_sig_loopback =3414;
22124: waveform_sig_loopback =1368;
22125: waveform_sig_loopback =3621;
22126: waveform_sig_loopback =2883;
22127: waveform_sig_loopback =1917;
22128: waveform_sig_loopback =2596;
22129: waveform_sig_loopback =3519;
22130: waveform_sig_loopback =1656;
22131: waveform_sig_loopback =1902;
22132: waveform_sig_loopback =3829;
22133: waveform_sig_loopback =1933;
22134: waveform_sig_loopback =1228;
22135: waveform_sig_loopback =3196;
22136: waveform_sig_loopback =2938;
22137: waveform_sig_loopback =1162;
22138: waveform_sig_loopback =1619;
22139: waveform_sig_loopback =3904;
22140: waveform_sig_loopback =939;
22141: waveform_sig_loopback =2880;
22142: waveform_sig_loopback =2090;
22143: waveform_sig_loopback =-1280;
22144: waveform_sig_loopback =4619;
22145: waveform_sig_loopback =2658;
22146: waveform_sig_loopback =529;
22147: waveform_sig_loopback =981;
22148: waveform_sig_loopback =1833;
22149: waveform_sig_loopback =3130;
22150: waveform_sig_loopback =1620;
22151: waveform_sig_loopback =85;
22152: waveform_sig_loopback =2454;
22153: waveform_sig_loopback =1265;
22154: waveform_sig_loopback =1776;
22155: waveform_sig_loopback =990;
22156: waveform_sig_loopback =1006;
22157: waveform_sig_loopback =2351;
22158: waveform_sig_loopback =435;
22159: waveform_sig_loopback =1372;
22160: waveform_sig_loopback =1146;
22161: waveform_sig_loopback =1417;
22162: waveform_sig_loopback =271;
22163: waveform_sig_loopback =1761;
22164: waveform_sig_loopback =1281;
22165: waveform_sig_loopback =-362;
22166: waveform_sig_loopback =1909;
22167: waveform_sig_loopback =957;
22168: waveform_sig_loopback =21;
22169: waveform_sig_loopback =892;
22170: waveform_sig_loopback =1644;
22171: waveform_sig_loopback =-299;
22172: waveform_sig_loopback =320;
22173: waveform_sig_loopback =1744;
22174: waveform_sig_loopback =129;
22175: waveform_sig_loopback =-552;
22176: waveform_sig_loopback =1139;
22177: waveform_sig_loopback =1331;
22178: waveform_sig_loopback =-1029;
22179: waveform_sig_loopback =-164;
22180: waveform_sig_loopback =2267;
22181: waveform_sig_loopback =-1454;
22182: waveform_sig_loopback =1543;
22183: waveform_sig_loopback =-178;
22184: waveform_sig_loopback =-3209;
22185: waveform_sig_loopback =3254;
22186: waveform_sig_loopback =192;
22187: waveform_sig_loopback =-1209;
22188: waveform_sig_loopback =-791;
22189: waveform_sig_loopback =-298;
22190: waveform_sig_loopback =1544;
22191: waveform_sig_loopback =-635;
22192: waveform_sig_loopback =-1793;
22193: waveform_sig_loopback =866;
22194: waveform_sig_loopback =-919;
22195: waveform_sig_loopback =45;
22196: waveform_sig_loopback =-893;
22197: waveform_sig_loopback =-1000;
22198: waveform_sig_loopback =657;
22199: waveform_sig_loopback =-1575;
22200: waveform_sig_loopback =-555;
22201: waveform_sig_loopback =-623;
22202: waveform_sig_loopback =-561;
22203: waveform_sig_loopback =-1690;
22204: waveform_sig_loopback =31;
22205: waveform_sig_loopback =-764;
22206: waveform_sig_loopback =-2248;
22207: waveform_sig_loopback =244;
22208: waveform_sig_loopback =-1255;
22209: waveform_sig_loopback =-1663;
22210: waveform_sig_loopback =-854;
22211: waveform_sig_loopback =-621;
22212: waveform_sig_loopback =-1829;
22213: waveform_sig_loopback =-1790;
22214: waveform_sig_loopback =-106;
22215: waveform_sig_loopback =-1606;
22216: waveform_sig_loopback =-2776;
22217: waveform_sig_loopback =-280;
22218: waveform_sig_loopback =-768;
22219: waveform_sig_loopback =-3114;
22220: waveform_sig_loopback =-1528;
22221: waveform_sig_loopback =9;
22222: waveform_sig_loopback =-3251;
22223: waveform_sig_loopback =-57;
22224: waveform_sig_loopback =-2606;
22225: waveform_sig_loopback =-4577;
22226: waveform_sig_loopback =1315;
22227: waveform_sig_loopback =-1926;
22228: waveform_sig_loopback =-2712;
22229: waveform_sig_loopback =-2940;
22230: waveform_sig_loopback =-2003;
22231: waveform_sig_loopback =-156;
22232: waveform_sig_loopback =-2801;
22233: waveform_sig_loopback =-3427;
22234: waveform_sig_loopback =-1068;
22235: waveform_sig_loopback =-2915;
22236: waveform_sig_loopback =-1611;
22237: waveform_sig_loopback =-2942;
22238: waveform_sig_loopback =-2797;
22239: waveform_sig_loopback =-1084;
22240: waveform_sig_loopback =-3580;
22241: waveform_sig_loopback =-2359;
22242: waveform_sig_loopback =-2309;
22243: waveform_sig_loopback =-2652;
22244: waveform_sig_loopback =-3353;
22245: waveform_sig_loopback =-1692;
22246: waveform_sig_loopback =-3017;
22247: waveform_sig_loopback =-3609;
22248: waveform_sig_loopback =-1871;
22249: waveform_sig_loopback =-3080;
22250: waveform_sig_loopback =-3262;
22251: waveform_sig_loopback =-3020;
22252: waveform_sig_loopback =-2045;
22253: waveform_sig_loopback =-3892;
22254: waveform_sig_loopback =-3590;
22255: waveform_sig_loopback =-1644;
22256: waveform_sig_loopback =-3751;
22257: waveform_sig_loopback =-4388;
22258: waveform_sig_loopback =-2009;
22259: waveform_sig_loopback =-2737;
22260: waveform_sig_loopback =-4812;
22261: waveform_sig_loopback =-3211;
22262: waveform_sig_loopback =-1942;
22263: waveform_sig_loopback =-4942;
22264: waveform_sig_loopback =-1680;
22265: waveform_sig_loopback =-4744;
22266: waveform_sig_loopback =-5945;
22267: waveform_sig_loopback =-505;
22268: waveform_sig_loopback =-3802;
22269: waveform_sig_loopback =-4277;
22270: waveform_sig_loopback =-4921;
22271: waveform_sig_loopback =-3434;
22272: waveform_sig_loopback =-1882;
22273: waveform_sig_loopback =-4849;
22274: waveform_sig_loopback =-4737;
22275: waveform_sig_loopback =-2986;
22276: waveform_sig_loopback =-4588;
22277: waveform_sig_loopback =-3096;
22278: waveform_sig_loopback =-5027;
22279: waveform_sig_loopback =-4063;
22280: waveform_sig_loopback =-2891;
22281: waveform_sig_loopback =-5407;
22282: waveform_sig_loopback =-3710;
22283: waveform_sig_loopback =-4189;
22284: waveform_sig_loopback =-4294;
22285: waveform_sig_loopback =-4862;
22286: waveform_sig_loopback =-3460;
22287: waveform_sig_loopback =-4648;
22288: waveform_sig_loopback =-5159;
22289: waveform_sig_loopback =-3644;
22290: waveform_sig_loopback =-4510;
22291: waveform_sig_loopback =-5018;
22292: waveform_sig_loopback =-4629;
22293: waveform_sig_loopback =-3461;
22294: waveform_sig_loopback =-5773;
22295: waveform_sig_loopback =-4996;
22296: waveform_sig_loopback =-3137;
22297: waveform_sig_loopback =-5579;
22298: waveform_sig_loopback =-5698;
22299: waveform_sig_loopback =-3631;
22300: waveform_sig_loopback =-4473;
22301: waveform_sig_loopback =-6100;
22302: waveform_sig_loopback =-4736;
22303: waveform_sig_loopback =-3661;
22304: waveform_sig_loopback =-6325;
22305: waveform_sig_loopback =-3148;
22306: waveform_sig_loopback =-6431;
22307: waveform_sig_loopback =-7228;
22308: waveform_sig_loopback =-2192;
22309: waveform_sig_loopback =-5076;
22310: waveform_sig_loopback =-5899;
22311: waveform_sig_loopback =-6565;
22312: waveform_sig_loopback =-4487;
22313: waveform_sig_loopback =-3655;
22314: waveform_sig_loopback =-6369;
22315: waveform_sig_loopback =-5981;
22316: waveform_sig_loopback =-4613;
22317: waveform_sig_loopback =-5758;
22318: waveform_sig_loopback =-4712;
22319: waveform_sig_loopback =-6527;
22320: waveform_sig_loopback =-5078;
22321: waveform_sig_loopback =-4654;
22322: waveform_sig_loopback =-6683;
22323: waveform_sig_loopback =-5034;
22324: waveform_sig_loopback =-5672;
22325: waveform_sig_loopback =-5494;
22326: waveform_sig_loopback =-6298;
22327: waveform_sig_loopback =-4791;
22328: waveform_sig_loopback =-6010;
22329: waveform_sig_loopback =-6414;
22330: waveform_sig_loopback =-5031;
22331: waveform_sig_loopback =-5811;
22332: waveform_sig_loopback =-6424;
22333: waveform_sig_loopback =-5840;
22334: waveform_sig_loopback =-4704;
22335: waveform_sig_loopback =-7377;
22336: waveform_sig_loopback =-5892;
22337: waveform_sig_loopback =-4459;
22338: waveform_sig_loopback =-7198;
22339: waveform_sig_loopback =-6583;
22340: waveform_sig_loopback =-4924;
22341: waveform_sig_loopback =-5728;
22342: waveform_sig_loopback =-7408;
22343: waveform_sig_loopback =-6051;
22344: waveform_sig_loopback =-4507;
22345: waveform_sig_loopback =-7655;
22346: waveform_sig_loopback =-4542;
22347: waveform_sig_loopback =-7495;
22348: waveform_sig_loopback =-8305;
22349: waveform_sig_loopback =-3275;
22350: waveform_sig_loopback =-6318;
22351: waveform_sig_loopback =-7208;
22352: waveform_sig_loopback =-7317;
22353: waveform_sig_loopback =-5751;
22354: waveform_sig_loopback =-4813;
22355: waveform_sig_loopback =-7180;
22356: waveform_sig_loopback =-7196;
22357: waveform_sig_loopback =-5689;
22358: waveform_sig_loopback =-6716;
22359: waveform_sig_loopback =-5802;
22360: waveform_sig_loopback =-7543;
22361: waveform_sig_loopback =-6024;
22362: waveform_sig_loopback =-5901;
22363: waveform_sig_loopback =-7444;
22364: waveform_sig_loopback =-6045;
22365: waveform_sig_loopback =-6820;
22366: waveform_sig_loopback =-6285;
22367: waveform_sig_loopback =-7379;
22368: waveform_sig_loopback =-5631;
22369: waveform_sig_loopback =-6893;
22370: waveform_sig_loopback =-7537;
22371: waveform_sig_loopback =-5624;
22372: waveform_sig_loopback =-6815;
22373: waveform_sig_loopback =-7559;
22374: waveform_sig_loopback =-6170;
22375: waveform_sig_loopback =-6006;
22376: waveform_sig_loopback =-8136;
22377: waveform_sig_loopback =-6487;
22378: waveform_sig_loopback =-5659;
22379: waveform_sig_loopback =-7676;
22380: waveform_sig_loopback =-7550;
22381: waveform_sig_loopback =-5752;
22382: waveform_sig_loopback =-6339;
22383: waveform_sig_loopback =-8416;
22384: waveform_sig_loopback =-6611;
22385: waveform_sig_loopback =-5299;
22386: waveform_sig_loopback =-8558;
22387: waveform_sig_loopback =-5014;
22388: waveform_sig_loopback =-8527;
22389: waveform_sig_loopback =-8922;
22390: waveform_sig_loopback =-3784;
22391: waveform_sig_loopback =-7221;
22392: waveform_sig_loopback =-8023;
22393: waveform_sig_loopback =-7714;
22394: waveform_sig_loopback =-6534;
22395: waveform_sig_loopback =-5502;
22396: waveform_sig_loopback =-7807;
22397: waveform_sig_loopback =-8039;
22398: waveform_sig_loopback =-6018;
22399: waveform_sig_loopback =-7480;
22400: waveform_sig_loopback =-6609;
22401: waveform_sig_loopback =-7784;
22402: waveform_sig_loopback =-6858;
22403: waveform_sig_loopback =-6408;
22404: waveform_sig_loopback =-7988;
22405: waveform_sig_loopback =-6776;
22406: waveform_sig_loopback =-7114;
22407: waveform_sig_loopback =-6962;
22408: waveform_sig_loopback =-8176;
22409: waveform_sig_loopback =-5848;
22410: waveform_sig_loopback =-7511;
22411: waveform_sig_loopback =-8024;
22412: waveform_sig_loopback =-6102;
22413: waveform_sig_loopback =-7546;
22414: waveform_sig_loopback =-7628;
22415: waveform_sig_loopback =-6583;
22416: waveform_sig_loopback =-6841;
22417: waveform_sig_loopback =-8259;
22418: waveform_sig_loopback =-6821;
22419: waveform_sig_loopback =-6190;
22420: waveform_sig_loopback =-8014;
22421: waveform_sig_loopback =-8112;
22422: waveform_sig_loopback =-5862;
22423: waveform_sig_loopback =-6784;
22424: waveform_sig_loopback =-9041;
22425: waveform_sig_loopback =-6513;
22426: waveform_sig_loopback =-5845;
22427: waveform_sig_loopback =-8921;
22428: waveform_sig_loopback =-5080;
22429: waveform_sig_loopback =-9281;
22430: waveform_sig_loopback =-8784;
22431: waveform_sig_loopback =-4029;
22432: waveform_sig_loopback =-7866;
22433: waveform_sig_loopback =-8018;
22434: waveform_sig_loopback =-8018;
22435: waveform_sig_loopback =-6885;
22436: waveform_sig_loopback =-5471;
22437: waveform_sig_loopback =-8323;
22438: waveform_sig_loopback =-8057;
22439: waveform_sig_loopback =-6060;
22440: waveform_sig_loopback =-7989;
22441: waveform_sig_loopback =-6385;
22442: waveform_sig_loopback =-8171;
22443: waveform_sig_loopback =-7029;
22444: waveform_sig_loopback =-6333;
22445: waveform_sig_loopback =-8303;
22446: waveform_sig_loopback =-6776;
22447: waveform_sig_loopback =-7094;
22448: waveform_sig_loopback =-7253;
22449: waveform_sig_loopback =-7819;
22450: waveform_sig_loopback =-5937;
22451: waveform_sig_loopback =-7889;
22452: waveform_sig_loopback =-7673;
22453: waveform_sig_loopback =-6033;
22454: waveform_sig_loopback =-7642;
22455: waveform_sig_loopback =-7588;
22456: waveform_sig_loopback =-6603;
22457: waveform_sig_loopback =-6645;
22458: waveform_sig_loopback =-8099;
22459: waveform_sig_loopback =-7084;
22460: waveform_sig_loopback =-5848;
22461: waveform_sig_loopback =-7881;
22462: waveform_sig_loopback =-8199;
22463: waveform_sig_loopback =-5395;
22464: waveform_sig_loopback =-6965;
22465: waveform_sig_loopback =-8811;
22466: waveform_sig_loopback =-5983;
22467: waveform_sig_loopback =-6255;
22468: waveform_sig_loopback =-8306;
22469: waveform_sig_loopback =-4839;
22470: waveform_sig_loopback =-9516;
22471: waveform_sig_loopback =-7910;
22472: waveform_sig_loopback =-4189;
22473: waveform_sig_loopback =-7495;
22474: waveform_sig_loopback =-7565;
22475: waveform_sig_loopback =-8149;
22476: waveform_sig_loopback =-6083;
22477: waveform_sig_loopback =-5225;
22478: waveform_sig_loopback =-8357;
22479: waveform_sig_loopback =-7363;
22480: waveform_sig_loopback =-5985;
22481: waveform_sig_loopback =-7468;
22482: waveform_sig_loopback =-5935;
22483: waveform_sig_loopback =-8065;
22484: waveform_sig_loopback =-6276;
22485: waveform_sig_loopback =-6033;
22486: waveform_sig_loopback =-7945;
22487: waveform_sig_loopback =-6184;
22488: waveform_sig_loopback =-6651;
22489: waveform_sig_loopback =-6922;
22490: waveform_sig_loopback =-7203;
22491: waveform_sig_loopback =-5508;
22492: waveform_sig_loopback =-7673;
22493: waveform_sig_loopback =-6761;
22494: waveform_sig_loopback =-5905;
22495: waveform_sig_loopback =-6947;
22496: waveform_sig_loopback =-6956;
22497: waveform_sig_loopback =-6435;
22498: waveform_sig_loopback =-5648;
22499: waveform_sig_loopback =-7929;
22500: waveform_sig_loopback =-6359;
22501: waveform_sig_loopback =-5025;
22502: waveform_sig_loopback =-7834;
22503: waveform_sig_loopback =-7072;
22504: waveform_sig_loopback =-4911;
22505: waveform_sig_loopback =-6584;
22506: waveform_sig_loopback =-7816;
22507: waveform_sig_loopback =-5589;
22508: waveform_sig_loopback =-5525;
22509: waveform_sig_loopback =-7499;
22510: waveform_sig_loopback =-4359;
22511: waveform_sig_loopback =-8848;
22512: waveform_sig_loopback =-7023;
22513: waveform_sig_loopback =-3574;
22514: waveform_sig_loopback =-6732;
22515: waveform_sig_loopback =-6940;
22516: waveform_sig_loopback =-7331;
22517: waveform_sig_loopback =-5160;
22518: waveform_sig_loopback =-4643;
22519: waveform_sig_loopback =-7637;
22520: waveform_sig_loopback =-6285;
22521: waveform_sig_loopback =-5419;
22522: waveform_sig_loopback =-6535;
22523: waveform_sig_loopback =-5039;
22524: waveform_sig_loopback =-7465;
22525: waveform_sig_loopback =-5055;
22526: waveform_sig_loopback =-5431;
22527: waveform_sig_loopback =-7127;
22528: waveform_sig_loopback =-5027;
22529: waveform_sig_loopback =-6126;
22530: waveform_sig_loopback =-5863;
22531: waveform_sig_loopback =-6092;
22532: waveform_sig_loopback =-4944;
22533: waveform_sig_loopback =-6330;
22534: waveform_sig_loopback =-6055;
22535: waveform_sig_loopback =-4994;
22536: waveform_sig_loopback =-5689;
22537: waveform_sig_loopback =-6458;
22538: waveform_sig_loopback =-4976;
22539: waveform_sig_loopback =-4885;
22540: waveform_sig_loopback =-7079;
22541: waveform_sig_loopback =-4958;
22542: waveform_sig_loopback =-4391;
22543: waveform_sig_loopback =-6755;
22544: waveform_sig_loopback =-5797;
22545: waveform_sig_loopback =-4022;
22546: waveform_sig_loopback =-5488;
22547: waveform_sig_loopback =-6689;
22548: waveform_sig_loopback =-4484;
22549: waveform_sig_loopback =-4425;
22550: waveform_sig_loopback =-6396;
22551: waveform_sig_loopback =-3304;
22552: waveform_sig_loopback =-7737;
22553: waveform_sig_loopback =-5694;
22554: waveform_sig_loopback =-2496;
22555: waveform_sig_loopback =-5538;
22556: waveform_sig_loopback =-5949;
22557: waveform_sig_loopback =-5996;
22558: waveform_sig_loopback =-3811;
22559: waveform_sig_loopback =-3785;
22560: waveform_sig_loopback =-6208;
22561: waveform_sig_loopback =-5026;
22562: waveform_sig_loopback =-4412;
22563: waveform_sig_loopback =-4952;
22564: waveform_sig_loopback =-4207;
22565: waveform_sig_loopback =-6034;
22566: waveform_sig_loopback =-3544;
22567: waveform_sig_loopback =-4674;
22568: waveform_sig_loopback =-5377;
22569: waveform_sig_loopback =-3909;
22570: waveform_sig_loopback =-4963;
22571: waveform_sig_loopback =-4211;
22572: waveform_sig_loopback =-5204;
22573: waveform_sig_loopback =-3272;
22574: waveform_sig_loopback =-5066;
22575: waveform_sig_loopback =-4940;
22576: waveform_sig_loopback =-3208;
22577: waveform_sig_loopback =-4733;
22578: waveform_sig_loopback =-4945;
22579: waveform_sig_loopback =-3418;
22580: waveform_sig_loopback =-3890;
22581: waveform_sig_loopback =-5385;
22582: waveform_sig_loopback =-3583;
22583: waveform_sig_loopback =-3020;
22584: waveform_sig_loopback =-5361;
22585: waveform_sig_loopback =-4310;
22586: waveform_sig_loopback =-2569;
22587: waveform_sig_loopback =-4199;
22588: waveform_sig_loopback =-5130;
22589: waveform_sig_loopback =-3123;
22590: waveform_sig_loopback =-2859;
22591: waveform_sig_loopback =-4962;
22592: waveform_sig_loopback =-1920;
22593: waveform_sig_loopback =-6105;
22594: waveform_sig_loopback =-4372;
22595: waveform_sig_loopback =-808;
22596: waveform_sig_loopback =-4083;
22597: waveform_sig_loopback =-4737;
22598: waveform_sig_loopback =-3960;
22599: waveform_sig_loopback =-2635;
22600: waveform_sig_loopback =-2166;
22601: waveform_sig_loopback =-4530;
22602: waveform_sig_loopback =-3855;
22603: waveform_sig_loopback =-2440;
22604: waveform_sig_loopback =-3579;
22605: waveform_sig_loopback =-2734;
22606: waveform_sig_loopback =-4117;
22607: waveform_sig_loopback =-2348;
22608: waveform_sig_loopback =-2904;
22609: waveform_sig_loopback =-3721;
22610: waveform_sig_loopback =-2620;
22611: waveform_sig_loopback =-2983;
22612: waveform_sig_loopback =-2889;
22613: waveform_sig_loopback =-3453;
22614: waveform_sig_loopback =-1587;
22615: waveform_sig_loopback =-3710;
22616: waveform_sig_loopback =-3031;
22617: waveform_sig_loopback =-1648;
22618: waveform_sig_loopback =-3107;
22619: waveform_sig_loopback =-3262;
22620: waveform_sig_loopback =-1604;
22621: waveform_sig_loopback =-2375;
22622: waveform_sig_loopback =-3634;
22623: waveform_sig_loopback =-1719;
22624: waveform_sig_loopback =-1659;
22625: waveform_sig_loopback =-3409;
22626: waveform_sig_loopback =-2721;
22627: waveform_sig_loopback =-892;
22628: waveform_sig_loopback =-2268;
22629: waveform_sig_loopback =-3798;
22630: waveform_sig_loopback =-954;
22631: waveform_sig_loopback =-1314;
22632: waveform_sig_loopback =-3404;
22633: waveform_sig_loopback =268;
22634: waveform_sig_loopback =-4960;
22635: waveform_sig_loopback =-2176;
22636: waveform_sig_loopback =1114;
22637: waveform_sig_loopback =-2889;
22638: waveform_sig_loopback =-2501;
22639: waveform_sig_loopback =-2336;
22640: waveform_sig_loopback =-940;
22641: waveform_sig_loopback =-83;
22642: waveform_sig_loopback =-3251;
22643: waveform_sig_loopback =-1676;
22644: waveform_sig_loopback =-688;
22645: waveform_sig_loopback =-2023;
22646: waveform_sig_loopback =-718;
22647: waveform_sig_loopback =-2446;
22648: waveform_sig_loopback =-497;
22649: waveform_sig_loopback =-1036;
22650: waveform_sig_loopback =-2021;
22651: waveform_sig_loopback =-726;
22652: waveform_sig_loopback =-1076;
22653: waveform_sig_loopback =-1235;
22654: waveform_sig_loopback =-1500;
22655: waveform_sig_loopback =352;
22656: waveform_sig_loopback =-2134;
22657: waveform_sig_loopback =-939;
22658: waveform_sig_loopback =114;
22659: waveform_sig_loopback =-1466;
22660: waveform_sig_loopback =-1157;
22661: waveform_sig_loopback =82;
22662: waveform_sig_loopback =-581;
22663: waveform_sig_loopback =-1651;
22664: waveform_sig_loopback =-46;
22665: waveform_sig_loopback =336;
22666: waveform_sig_loopback =-1570;
22667: waveform_sig_loopback =-961;
22668: waveform_sig_loopback =1242;
22669: waveform_sig_loopback =-678;
22670: waveform_sig_loopback =-1937;
22671: waveform_sig_loopback =1328;
22672: waveform_sig_loopback =-35;
22673: waveform_sig_loopback =-1123;
22674: waveform_sig_loopback =2158;
22675: waveform_sig_loopback =-3586;
22676: waveform_sig_loopback =471;
22677: waveform_sig_loopback =2458;
22678: waveform_sig_loopback =-932;
22679: waveform_sig_loopback =-381;
22680: waveform_sig_loopback =-897;
22681: waveform_sig_loopback =1454;
22682: waveform_sig_loopback =1519;
22683: waveform_sig_loopback =-1547;
22684: waveform_sig_loopback =601;
22685: waveform_sig_loopback =826;
22686: waveform_sig_loopback =71;
22687: waveform_sig_loopback =1105;
22688: waveform_sig_loopback =-760;
22689: waveform_sig_loopback =1638;
22690: waveform_sig_loopback =671;
22691: waveform_sig_loopback =-119;
22692: waveform_sig_loopback =1146;
22693: waveform_sig_loopback =884;
22694: waveform_sig_loopback =459;
22695: waveform_sig_loopback =580;
22696: waveform_sig_loopback =2111;
22697: waveform_sig_loopback =-490;
22698: waveform_sig_loopback =1418;
22699: waveform_sig_loopback =1604;
22700: waveform_sig_loopback =562;
22701: waveform_sig_loopback =858;
22702: waveform_sig_loopback =1582;
22703: waveform_sig_loopback =1772;
22704: waveform_sig_loopback =-80;
22705: waveform_sig_loopback =1978;
22706: waveform_sig_loopback =2373;
22707: waveform_sig_loopback =-123;
22708: waveform_sig_loopback =1446;
22709: waveform_sig_loopback =2916;
22710: waveform_sig_loopback =981;
22711: waveform_sig_loopback =264;
22712: waveform_sig_loopback =3122;
22713: waveform_sig_loopback =1736;
22714: waveform_sig_loopback =1042;
22715: waveform_sig_loopback =3765;
22716: waveform_sig_loopback =-1752;
22717: waveform_sig_loopback =2742;
22718: waveform_sig_loopback =3981;
22719: waveform_sig_loopback =1169;
22720: waveform_sig_loopback =1349;
22721: waveform_sig_loopback =926;
22722: waveform_sig_loopback =3725;
22723: waveform_sig_loopback =3016;
22724: waveform_sig_loopback =424;
22725: waveform_sig_loopback =2676;
22726: waveform_sig_loopback =2392;
22727: waveform_sig_loopback =2278;
22728: waveform_sig_loopback =2848;
22729: waveform_sig_loopback =1039;
22730: waveform_sig_loopback =3798;
22731: waveform_sig_loopback =2268;
22732: waveform_sig_loopback =1867;
22733: waveform_sig_loopback =3130;
22734: waveform_sig_loopback =2559;
22735: waveform_sig_loopback =2367;
22736: waveform_sig_loopback =2582;
22737: waveform_sig_loopback =3741;
22738: waveform_sig_loopback =1541;
22739: waveform_sig_loopback =3240;
22740: waveform_sig_loopback =3267;
22741: waveform_sig_loopback =2660;
22742: waveform_sig_loopback =2454;
22743: waveform_sig_loopback =3647;
22744: waveform_sig_loopback =3495;
22745: waveform_sig_loopback =1470;
22746: waveform_sig_loopback =4178;
22747: waveform_sig_loopback =3985;
22748: waveform_sig_loopback =1497;
22749: waveform_sig_loopback =3573;
22750: waveform_sig_loopback =4516;
22751: waveform_sig_loopback =2708;
22752: waveform_sig_loopback =2188;
22753: waveform_sig_loopback =4669;
22754: waveform_sig_loopback =3608;
22755: waveform_sig_loopback =2862;
22756: waveform_sig_loopback =5096;
22757: waveform_sig_loopback =178;
22758: waveform_sig_loopback =4541;
22759: waveform_sig_loopback =5697;
22760: waveform_sig_loopback =2817;
22761: waveform_sig_loopback =2606;
22762: waveform_sig_loopback =3245;
22763: waveform_sig_loopback =5368;
22764: waveform_sig_loopback =4429;
22765: waveform_sig_loopback =2220;
22766: waveform_sig_loopback =4417;
22767: waveform_sig_loopback =4159;
22768: waveform_sig_loopback =3893;
22769: waveform_sig_loopback =4324;
22770: waveform_sig_loopback =2904;
22771: waveform_sig_loopback =5554;
22772: waveform_sig_loopback =3610;
22773: waveform_sig_loopback =3679;
22774: waveform_sig_loopback =4857;
22775: waveform_sig_loopback =4007;
22776: waveform_sig_loopback =4121;
22777: waveform_sig_loopback =4152;
22778: waveform_sig_loopback =5315;
22779: waveform_sig_loopback =3416;
22780: waveform_sig_loopback =4464;
22781: waveform_sig_loopback =5144;
22782: waveform_sig_loopback =4254;
22783: waveform_sig_loopback =3728;
22784: waveform_sig_loopback =5712;
22785: waveform_sig_loopback =4559;
22786: waveform_sig_loopback =3271;
22787: waveform_sig_loopback =5994;
22788: waveform_sig_loopback =5009;
22789: waveform_sig_loopback =3430;
22790: waveform_sig_loopback =5067;
22791: waveform_sig_loopback =5958;
22792: waveform_sig_loopback =4400;
22793: waveform_sig_loopback =3579;
22794: waveform_sig_loopback =6431;
22795: waveform_sig_loopback =5039;
22796: waveform_sig_loopback =4299;
22797: waveform_sig_loopback =6825;
22798: waveform_sig_loopback =1610;
22799: waveform_sig_loopback =6005;
22800: waveform_sig_loopback =7249;
22801: waveform_sig_loopback =4236;
22802: waveform_sig_loopback =4218;
22803: waveform_sig_loopback =4723;
22804: waveform_sig_loopback =6599;
22805: waveform_sig_loopback =5996;
22806: waveform_sig_loopback =3851;
22807: waveform_sig_loopback =5632;
22808: waveform_sig_loopback =5594;
22809: waveform_sig_loopback =5449;
22810: waveform_sig_loopback =5542;
22811: waveform_sig_loopback =4532;
22812: waveform_sig_loopback =6738;
22813: waveform_sig_loopback =4958;
22814: waveform_sig_loopback =5382;
22815: waveform_sig_loopback =5868;
22816: waveform_sig_loopback =5553;
22817: waveform_sig_loopback =5543;
22818: waveform_sig_loopback =5280;
22819: waveform_sig_loopback =6904;
22820: waveform_sig_loopback =4439;
22821: waveform_sig_loopback =5908;
22822: waveform_sig_loopback =6689;
22823: waveform_sig_loopback =4989;
22824: waveform_sig_loopback =5433;
22825: waveform_sig_loopback =7021;
22826: waveform_sig_loopback =5448;
22827: waveform_sig_loopback =4948;
22828: waveform_sig_loopback =6964;
22829: waveform_sig_loopback =6283;
22830: waveform_sig_loopback =4798;
22831: waveform_sig_loopback =6028;
22832: waveform_sig_loopback =7401;
22833: waveform_sig_loopback =5422;
22834: waveform_sig_loopback =4749;
22835: waveform_sig_loopback =7891;
22836: waveform_sig_loopback =5870;
22837: waveform_sig_loopback =5703;
22838: waveform_sig_loopback =7892;
22839: waveform_sig_loopback =2653;
22840: waveform_sig_loopback =7482;
22841: waveform_sig_loopback =8191;
22842: waveform_sig_loopback =5310;
22843: waveform_sig_loopback =5346;
22844: waveform_sig_loopback =5913;
22845: waveform_sig_loopback =7598;
22846: waveform_sig_loopback =7115;
22847: waveform_sig_loopback =4852;
22848: waveform_sig_loopback =6584;
22849: waveform_sig_loopback =6893;
22850: waveform_sig_loopback =6291;
22851: waveform_sig_loopback =6593;
22852: waveform_sig_loopback =5744;
22853: waveform_sig_loopback =7476;
22854: waveform_sig_loopback =6275;
22855: waveform_sig_loopback =6205;
22856: waveform_sig_loopback =6665;
22857: waveform_sig_loopback =6976;
22858: waveform_sig_loopback =5979;
22859: waveform_sig_loopback =6629;
22860: waveform_sig_loopback =7802;
22861: waveform_sig_loopback =4995;
22862: waveform_sig_loopback =7461;
22863: waveform_sig_loopback =7117;
22864: waveform_sig_loopback =6071;
22865: waveform_sig_loopback =6499;
22866: waveform_sig_loopback =7607;
22867: waveform_sig_loopback =6613;
22868: waveform_sig_loopback =5652;
22869: waveform_sig_loopback =7920;
22870: waveform_sig_loopback =7118;
22871: waveform_sig_loopback =5519;
22872: waveform_sig_loopback =6997;
22873: waveform_sig_loopback =8165;
22874: waveform_sig_loopback =6221;
22875: waveform_sig_loopback =5457;
22876: waveform_sig_loopback =8895;
22877: waveform_sig_loopback =6382;
22878: waveform_sig_loopback =6612;
22879: waveform_sig_loopback =8698;
22880: waveform_sig_loopback =2981;
22881: waveform_sig_loopback =8761;
22882: waveform_sig_loopback =8721;
22883: waveform_sig_loopback =5708;
22884: waveform_sig_loopback =6485;
22885: waveform_sig_loopback =6296;
22886: waveform_sig_loopback =8467;
22887: waveform_sig_loopback =7889;
22888: waveform_sig_loopback =5045;
22889: waveform_sig_loopback =7813;
22890: waveform_sig_loopback =7184;
22891: waveform_sig_loopback =6839;
22892: waveform_sig_loopback =7531;
22893: waveform_sig_loopback =5896;
22894: waveform_sig_loopback =8384;
22895: waveform_sig_loopback =6770;
22896: waveform_sig_loopback =6544;
22897: waveform_sig_loopback =7633;
22898: waveform_sig_loopback =7192;
22899: waveform_sig_loopback =6530;
22900: waveform_sig_loopback =7380;
22901: waveform_sig_loopback =7975;
22902: waveform_sig_loopback =5758;
22903: waveform_sig_loopback =7862;
22904: waveform_sig_loopback =7521;
22905: waveform_sig_loopback =6578;
22906: waveform_sig_loopback =6982;
22907: waveform_sig_loopback =8009;
22908: waveform_sig_loopback =6937;
22909: waveform_sig_loopback =6199;
22910: waveform_sig_loopback =8205;
22911: waveform_sig_loopback =7651;
22912: waveform_sig_loopback =5731;
22913: waveform_sig_loopback =7434;
22914: waveform_sig_loopback =8714;
22915: waveform_sig_loopback =6117;
22916: waveform_sig_loopback =6192;
22917: waveform_sig_loopback =9186;
22918: waveform_sig_loopback =6299;
22919: waveform_sig_loopback =7494;
22920: waveform_sig_loopback =8411;
22921: waveform_sig_loopback =3391;
22922: waveform_sig_loopback =9420;
22923: waveform_sig_loopback =8413;
22924: waveform_sig_loopback =6371;
22925: waveform_sig_loopback =6483;
22926: waveform_sig_loopback =6409;
22927: waveform_sig_loopback =9114;
22928: waveform_sig_loopback =7524;
22929: waveform_sig_loopback =5445;
22930: waveform_sig_loopback =8145;
22931: waveform_sig_loopback =6914;
22932: waveform_sig_loopback =7449;
22933: waveform_sig_loopback =7328;
22934: waveform_sig_loopback =6010;
22935: waveform_sig_loopback =8790;
22936: waveform_sig_loopback =6409;
22937: waveform_sig_loopback =6940;
22938: waveform_sig_loopback =7617;
22939: waveform_sig_loopback =7107;
22940: waveform_sig_loopback =6730;
22941: waveform_sig_loopback =7404;
22942: waveform_sig_loopback =7881;
22943: waveform_sig_loopback =5767;
22944: waveform_sig_loopback =7921;
22945: waveform_sig_loopback =7355;
22946: waveform_sig_loopback =6618;
22947: waveform_sig_loopback =6886;
22948: waveform_sig_loopback =7861;
22949: waveform_sig_loopback =7011;
22950: waveform_sig_loopback =5878;
22951: waveform_sig_loopback =8348;
22952: waveform_sig_loopback =7551;
22953: waveform_sig_loopback =5239;
22954: waveform_sig_loopback =7894;
22955: waveform_sig_loopback =8231;
22956: waveform_sig_loopback =5854;
22957: waveform_sig_loopback =6489;
22958: waveform_sig_loopback =8473;
22959: waveform_sig_loopback =6480;
22960: waveform_sig_loopback =7278;
22961: waveform_sig_loopback =7833;
22962: waveform_sig_loopback =3636;
22963: waveform_sig_loopback =8906;
22964: waveform_sig_loopback =8305;
22965: waveform_sig_loopback =6211;
22966: waveform_sig_loopback =5821;
22967: waveform_sig_loopback =6570;
22968: waveform_sig_loopback =8614;
22969: waveform_sig_loopback =7197;
22970: waveform_sig_loopback =5284;
22971: waveform_sig_loopback =7651;
22972: waveform_sig_loopback =6665;
22973: waveform_sig_loopback =7233;
22974: waveform_sig_loopback =6795;
22975: waveform_sig_loopback =5759;
22976: waveform_sig_loopback =8462;
22977: waveform_sig_loopback =5895;
22978: waveform_sig_loopback =6654;
22979: waveform_sig_loopback =7235;
22980: waveform_sig_loopback =6494;
22981: waveform_sig_loopback =6515;
22982: waveform_sig_loopback =6904;
22983: waveform_sig_loopback =7200;
22984: waveform_sig_loopback =5682;
22985: waveform_sig_loopback =7060;
22986: waveform_sig_loopback =7132;
22987: waveform_sig_loopback =6092;
22988: waveform_sig_loopback =6118;
22989: waveform_sig_loopback =7869;
22990: waveform_sig_loopback =5955;
22991: waveform_sig_loopback =5521;
22992: waveform_sig_loopback =7977;
22993: waveform_sig_loopback =6497;
22994: waveform_sig_loopback =5059;
22995: waveform_sig_loopback =7155;
22996: waveform_sig_loopback =7488;
22997: waveform_sig_loopback =5410;
22998: waveform_sig_loopback =5653;
22999: waveform_sig_loopback =8001;
23000: waveform_sig_loopback =5745;
23001: waveform_sig_loopback =6637;
23002: waveform_sig_loopback =7065;
23003: waveform_sig_loopback =2977;
23004: waveform_sig_loopback =8278;
23005: waveform_sig_loopback =7533;
23006: waveform_sig_loopback =5291;
23007: waveform_sig_loopback =5091;
23008: waveform_sig_loopback =6058;
23009: waveform_sig_loopback =7686;
23010: waveform_sig_loopback =6287;
23011: waveform_sig_loopback =4671;
23012: waveform_sig_loopback =6760;
23013: waveform_sig_loopback =5886;
23014: waveform_sig_loopback =6415;
23015: waveform_sig_loopback =5722;
23016: waveform_sig_loopback =5323;
23017: waveform_sig_loopback =7393;
23018: waveform_sig_loopback =4876;
23019: waveform_sig_loopback =6128;
23020: waveform_sig_loopback =5975;
23021: waveform_sig_loopback =5830;
23022: waveform_sig_loopback =5555;
23023: waveform_sig_loopback =5834;
23024: waveform_sig_loopback =6586;
23025: waveform_sig_loopback =4437;
23026: waveform_sig_loopback =6239;
23027: waveform_sig_loopback =6302;
23028: waveform_sig_loopback =4764;
23029: waveform_sig_loopback =5526;
23030: waveform_sig_loopback =6760;
23031: waveform_sig_loopback =4722;
23032: waveform_sig_loopback =4916;
23033: waveform_sig_loopback =6785;
23034: waveform_sig_loopback =5398;
23035: waveform_sig_loopback =4142;
23036: waveform_sig_loopback =6070;
23037: waveform_sig_loopback =6451;
23038: waveform_sig_loopback =4288;
23039: waveform_sig_loopback =4552;
23040: waveform_sig_loopback =7081;
23041: waveform_sig_loopback =4441;
23042: waveform_sig_loopback =5611;
23043: waveform_sig_loopback =5946;
23044: waveform_sig_loopback =1762;
23045: waveform_sig_loopback =7295;
23046: waveform_sig_loopback =6394;
23047: waveform_sig_loopback =3965;
23048: waveform_sig_loopback =4119;
23049: waveform_sig_loopback =4960;
23050: waveform_sig_loopback =6337;
23051: waveform_sig_loopback =5240;
23052: waveform_sig_loopback =3420;
23053: waveform_sig_loopback =5520;
23054: waveform_sig_loopback =4889;
23055: waveform_sig_loopback =4919;
23056: waveform_sig_loopback =4628;
23057: waveform_sig_loopback =4199;
23058: waveform_sig_loopback =5801;
23059: waveform_sig_loopback =3972;
23060: waveform_sig_loopback =4658;
23061: waveform_sig_loopback =4720;
23062: waveform_sig_loopback =4825;
23063: waveform_sig_loopback =3838;
23064: waveform_sig_loopback =4950;
23065: waveform_sig_loopback =5120;
23066: waveform_sig_loopback =2945;
23067: waveform_sig_loopback =5258;
23068: waveform_sig_loopback =4702;
23069: waveform_sig_loopback =3490;
23070: waveform_sig_loopback =4245;
23071: waveform_sig_loopback =5226;
23072: waveform_sig_loopback =3442;
23073: waveform_sig_loopback =3574;
23074: waveform_sig_loopback =5295;
23075: waveform_sig_loopback =3981;
23076: waveform_sig_loopback =2845;
23077: waveform_sig_loopback =4584;
23078: waveform_sig_loopback =5081;
23079: waveform_sig_loopback =2771;
23080: waveform_sig_loopback =3086;
23081: waveform_sig_loopback =5932;
23082: waveform_sig_loopback =2592;
23083: waveform_sig_loopback =4436;
23084: waveform_sig_loopback =4391;
23085: waveform_sig_loopback =5;
23086: waveform_sig_loopback =6424;
23087: waveform_sig_loopback =4515;
23088: waveform_sig_loopback =2334;
23089: waveform_sig_loopback =2954;
23090: waveform_sig_loopback =3077;
23091: waveform_sig_loopback =5125;
23092: waveform_sig_loopback =3606;
23093: waveform_sig_loopback =1547;
23094: waveform_sig_loopback =4442;
23095: waveform_sig_loopback =2985;
23096: waveform_sig_loopback =3488;
23097: waveform_sig_loopback =3120;
23098: waveform_sig_loopback =2431;
23099: waveform_sig_loopback =4377;
23100: waveform_sig_loopback =2310;
23101: waveform_sig_loopback =2929;
23102: waveform_sig_loopback =3263;
23103: waveform_sig_loopback =2940;
23104: waveform_sig_loopback =2136;
23105: waveform_sig_loopback =3637;
23106: waveform_sig_loopback =3250;
23107: waveform_sig_loopback =1212;
23108: waveform_sig_loopback =3706;
23109: waveform_sig_loopback =2994;
23110: waveform_sig_loopback =1870;
23111: waveform_sig_loopback =2700;
23112: waveform_sig_loopback =3200;
23113: waveform_sig_loopback =2073;
23114: waveform_sig_loopback =1912;
23115: waveform_sig_loopback =3361;
23116: waveform_sig_loopback =2510;
23117: waveform_sig_loopback =827;
23118: waveform_sig_loopback =3167;
23119: waveform_sig_loopback =3306;
23120: waveform_sig_loopback =651;
23121: waveform_sig_loopback =1958;
23122: waveform_sig_loopback =3890;
23123: waveform_sig_loopback =650;
23124: waveform_sig_loopback =3186;
23125: waveform_sig_loopback =2140;
23126: waveform_sig_loopback =-1423;
23127: waveform_sig_loopback =4737;
23128: waveform_sig_loopback =2362;
23129: waveform_sig_loopback =945;
23130: waveform_sig_loopback =939;
23131: waveform_sig_loopback =1291;
23132: waveform_sig_loopback =3700;
23133: waveform_sig_loopback =1420;
23134: waveform_sig_loopback =-78;
23135: waveform_sig_loopback =2723;
23136: waveform_sig_loopback =922;
23137: waveform_sig_loopback =2041;
23138: waveform_sig_loopback =1036;
23139: waveform_sig_loopback =615;
23140: waveform_sig_loopback =2866;
23141: waveform_sig_loopback =221;
23142: waveform_sig_loopback =1268;
23143: waveform_sig_loopback =1419;
23144: waveform_sig_loopback =1176;
23145: waveform_sig_loopback =399;
23146: waveform_sig_loopback =1778;
23147: waveform_sig_loopback =1121;
23148: waveform_sig_loopback =-209;
23149: waveform_sig_loopback =1962;
23150: waveform_sig_loopback =690;
23151: waveform_sig_loopback =338;
23152: waveform_sig_loopback =706;
23153: waveform_sig_loopback =1564;
23154: waveform_sig_loopback =121;
23155: waveform_sig_loopback =-249;
23156: waveform_sig_loopback =2036;
23157: waveform_sig_loopback =399;
23158: waveform_sig_loopback =-1122;
23159: waveform_sig_loopback =1640;
23160: waveform_sig_loopback =1208;
23161: waveform_sig_loopback =-1132;
23162: waveform_sig_loopback =207;
23163: waveform_sig_loopback =1793;
23164: waveform_sig_loopback =-956;
23165: waveform_sig_loopback =1393;
23166: waveform_sig_loopback =-274;
23167: waveform_sig_loopback =-2827;
23168: waveform_sig_loopback =2766;
23169: waveform_sig_loopback =402;
23170: waveform_sig_loopback =-773;
23171: waveform_sig_loopback =-1235;
23172: waveform_sig_loopback =-209;
23173: waveform_sig_loopback =1735;
23174: waveform_sig_loopback =-785;
23175: waveform_sig_loopback =-1610;
23176: waveform_sig_loopback =691;
23177: waveform_sig_loopback =-1037;
23178: waveform_sig_loopback =364;
23179: waveform_sig_loopback =-1176;
23180: waveform_sig_loopback =-998;
23181: waveform_sig_loopback =910;
23182: waveform_sig_loopback =-1920;
23183: waveform_sig_loopback =-349;
23184: waveform_sig_loopback =-602;
23185: waveform_sig_loopback =-860;
23186: waveform_sig_loopback =-1306;
23187: waveform_sig_loopback =-206;
23188: waveform_sig_loopback =-900;
23189: waveform_sig_loopback =-1881;
23190: waveform_sig_loopback =-216;
23191: waveform_sig_loopback =-1012;
23192: waveform_sig_loopback =-1581;
23193: waveform_sig_loopback =-1386;
23194: waveform_sig_loopback =24;
23195: waveform_sig_loopback =-2167;
23196: waveform_sig_loopback =-1986;
23197: waveform_sig_loopback =356;
23198: waveform_sig_loopback =-1972;
23199: waveform_sig_loopback =-2662;
23200: waveform_sig_loopback =-298;
23201: waveform_sig_loopback =-894;
23202: waveform_sig_loopback =-2819;
23203: waveform_sig_loopback =-1785;
23204: waveform_sig_loopback =-29;
23205: waveform_sig_loopback =-2805;
23206: waveform_sig_loopback =-475;
23207: waveform_sig_loopback =-2283;
23208: waveform_sig_loopback =-4483;
23209: waveform_sig_loopback =862;
23210: waveform_sig_loopback =-1481;
23211: waveform_sig_loopback =-2724;
23212: waveform_sig_loopback =-3193;
23213: waveform_sig_loopback =-1691;
23214: waveform_sig_loopback =-418;
23215: waveform_sig_loopback =-2670;
23216: waveform_sig_loopback =-3223;
23217: waveform_sig_loopback =-1428;
23218: waveform_sig_loopback =-2627;
23219: waveform_sig_loopback =-1630;
23220: waveform_sig_loopback =-3155;
23221: waveform_sig_loopback =-2483;
23222: waveform_sig_loopback =-1281;
23223: waveform_sig_loopback =-3669;
23224: waveform_sig_loopback =-2069;
23225: waveform_sig_loopback =-2561;
23226: waveform_sig_loopback =-2594;
23227: waveform_sig_loopback =-3204;
23228: waveform_sig_loopback =-2043;
23229: waveform_sig_loopback =-2661;
23230: waveform_sig_loopback =-3700;
23231: waveform_sig_loopback =-2101;
23232: waveform_sig_loopback =-2632;
23233: waveform_sig_loopback =-3607;
23234: waveform_sig_loopback =-3032;
23235: waveform_sig_loopback =-1678;
23236: waveform_sig_loopback =-4351;
23237: waveform_sig_loopback =-3320;
23238: waveform_sig_loopback =-1596;
23239: waveform_sig_loopback =-4022;
23240: waveform_sig_loopback =-3994;
23241: waveform_sig_loopback =-2410;
23242: waveform_sig_loopback =-2597;
23243: waveform_sig_loopback =-4541;
23244: waveform_sig_loopback =-3787;
23245: waveform_sig_loopback =-1498;
23246: waveform_sig_loopback =-4966;
23247: waveform_sig_loopback =-2096;
23248: waveform_sig_loopback =-4126;
23249: waveform_sig_loopback =-6367;
23250: waveform_sig_loopback =-580;
23251: waveform_sig_loopback =-3439;
23252: waveform_sig_loopback =-4620;
23253: waveform_sig_loopback =-4727;
23254: waveform_sig_loopback =-3451;
23255: waveform_sig_loopback =-2217;
23256: waveform_sig_loopback =-4398;
23257: waveform_sig_loopback =-4908;
23258: waveform_sig_loopback =-3130;
23259: waveform_sig_loopback =-4228;
23260: waveform_sig_loopback =-3511;
23261: waveform_sig_loopback =-4803;
23262: waveform_sig_loopback =-3975;
23263: waveform_sig_loopback =-3247;
23264: waveform_sig_loopback =-5132;
23265: waveform_sig_loopback =-3792;
23266: waveform_sig_loopback =-4391;
23267: waveform_sig_loopback =-3950;
23268: waveform_sig_loopback =-5092;
23269: waveform_sig_loopback =-3543;
23270: waveform_sig_loopback =-4227;
23271: waveform_sig_loopback =-5583;
23272: waveform_sig_loopback =-3391;
23273: waveform_sig_loopback =-4412;
23274: waveform_sig_loopback =-5410;
23275: waveform_sig_loopback =-4158;
23276: waveform_sig_loopback =-3776;
23277: waveform_sig_loopback =-5754;
23278: waveform_sig_loopback =-4732;
23279: waveform_sig_loopback =-3530;
23280: waveform_sig_loopback =-5326;
23281: waveform_sig_loopback =-5741;
23282: waveform_sig_loopback =-3836;
23283: waveform_sig_loopback =-4070;
23284: waveform_sig_loopback =-6371;
23285: waveform_sig_loopback =-4963;
23286: waveform_sig_loopback =-3107;
23287: waveform_sig_loopback =-6651;
23288: waveform_sig_loopback =-3352;
23289: waveform_sig_loopback =-5905;
23290: waveform_sig_loopback =-7736;
23291: waveform_sig_loopback =-1922;
23292: waveform_sig_loopback =-5099;
23293: waveform_sig_loopback =-6127;
23294: waveform_sig_loopback =-6040;
23295: waveform_sig_loopback =-4937;
23296: waveform_sig_loopback =-3667;
23297: waveform_sig_loopback =-5848;
23298: waveform_sig_loopback =-6510;
23299: waveform_sig_loopback =-4400;
23300: waveform_sig_loopback =-5644;
23301: waveform_sig_loopback =-5074;
23302: waveform_sig_loopback =-5989;
23303: waveform_sig_loopback =-5490;
23304: waveform_sig_loopback =-4643;
23305: waveform_sig_loopback =-6258;
23306: waveform_sig_loopback =-5488;
23307: waveform_sig_loopback =-5479;
23308: waveform_sig_loopback =-5317;
23309: waveform_sig_loopback =-6716;
23310: waveform_sig_loopback =-4430;
23311: waveform_sig_loopback =-6028;
23312: waveform_sig_loopback =-6777;
23313: waveform_sig_loopback =-4482;
23314: waveform_sig_loopback =-6200;
23315: waveform_sig_loopback =-6330;
23316: waveform_sig_loopback =-5615;
23317: waveform_sig_loopback =-5140;
23318: waveform_sig_loopback =-6848;
23319: waveform_sig_loopback =-6225;
23320: waveform_sig_loopback =-4595;
23321: waveform_sig_loopback =-6652;
23322: waveform_sig_loopback =-7050;
23323: waveform_sig_loopback =-4851;
23324: waveform_sig_loopback =-5458;
23325: waveform_sig_loopback =-7618;
23326: waveform_sig_loopback =-6010;
23327: waveform_sig_loopback =-4395;
23328: waveform_sig_loopback =-7882;
23329: waveform_sig_loopback =-4336;
23330: waveform_sig_loopback =-7406;
23331: waveform_sig_loopback =-8709;
23332: waveform_sig_loopback =-2857;
23333: waveform_sig_loopback =-6574;
23334: waveform_sig_loopback =-7176;
23335: waveform_sig_loopback =-7003;
23336: waveform_sig_loopback =-6312;
23337: waveform_sig_loopback =-4397;
23338: waveform_sig_loopback =-7249;
23339: waveform_sig_loopback =-7600;
23340: waveform_sig_loopback =-5093;
23341: waveform_sig_loopback =-7257;
23342: waveform_sig_loopback =-5707;
23343: waveform_sig_loopback =-7175;
23344: waveform_sig_loopback =-6725;
23345: waveform_sig_loopback =-5265;
23346: waveform_sig_loopback =-7747;
23347: waveform_sig_loopback =-6283;
23348: waveform_sig_loopback =-6341;
23349: waveform_sig_loopback =-6769;
23350: waveform_sig_loopback =-7185;
23351: waveform_sig_loopback =-5596;
23352: waveform_sig_loopback =-7104;
23353: waveform_sig_loopback =-7328;
23354: waveform_sig_loopback =-5767;
23355: waveform_sig_loopback =-6863;
23356: waveform_sig_loopback =-7347;
23357: waveform_sig_loopback =-6482;
23358: waveform_sig_loopback =-5961;
23359: waveform_sig_loopback =-7826;
23360: waveform_sig_loopback =-6913;
23361: waveform_sig_loopback =-5593;
23362: waveform_sig_loopback =-7379;
23363: waveform_sig_loopback =-8028;
23364: waveform_sig_loopback =-5482;
23365: waveform_sig_loopback =-6291;
23366: waveform_sig_loopback =-8671;
23367: waveform_sig_loopback =-6318;
23368: waveform_sig_loopback =-5663;
23369: waveform_sig_loopback =-8512;
23370: waveform_sig_loopback =-4759;
23371: waveform_sig_loopback =-8843;
23372: waveform_sig_loopback =-8694;
23373: waveform_sig_loopback =-3845;
23374: waveform_sig_loopback =-7508;
23375: waveform_sig_loopback =-7447;
23376: waveform_sig_loopback =-8283;
23377: waveform_sig_loopback =-6481;
23378: waveform_sig_loopback =-5115;
23379: waveform_sig_loopback =-8352;
23380: waveform_sig_loopback =-7629;
23381: waveform_sig_loopback =-6151;
23382: waveform_sig_loopback =-7751;
23383: waveform_sig_loopback =-6123;
23384: waveform_sig_loopback =-8228;
23385: waveform_sig_loopback =-6805;
23386: waveform_sig_loopback =-6068;
23387: waveform_sig_loopback =-8422;
23388: waveform_sig_loopback =-6511;
23389: waveform_sig_loopback =-7148;
23390: waveform_sig_loopback =-7167;
23391: waveform_sig_loopback =-7715;
23392: waveform_sig_loopback =-6111;
23393: waveform_sig_loopback =-7657;
23394: waveform_sig_loopback =-7745;
23395: waveform_sig_loopback =-6245;
23396: waveform_sig_loopback =-7387;
23397: waveform_sig_loopback =-7618;
23398: waveform_sig_loopback =-7050;
23399: waveform_sig_loopback =-6330;
23400: waveform_sig_loopback =-8204;
23401: waveform_sig_loopback =-7414;
23402: waveform_sig_loopback =-5640;
23403: waveform_sig_loopback =-8224;
23404: waveform_sig_loopback =-8178;
23405: waveform_sig_loopback =-5563;
23406: waveform_sig_loopback =-7212;
23407: waveform_sig_loopback =-8547;
23408: waveform_sig_loopback =-6712;
23409: waveform_sig_loopback =-6099;
23410: waveform_sig_loopback =-8380;
23411: waveform_sig_loopback =-5487;
23412: waveform_sig_loopback =-9009;
23413: waveform_sig_loopback =-8675;
23414: waveform_sig_loopback =-4466;
23415: waveform_sig_loopback =-7312;
23416: waveform_sig_loopback =-7923;
23417: waveform_sig_loopback =-8505;
23418: waveform_sig_loopback =-6338;
23419: waveform_sig_loopback =-5736;
23420: waveform_sig_loopback =-8273;
23421: waveform_sig_loopback =-7733;
23422: waveform_sig_loopback =-6614;
23423: waveform_sig_loopback =-7522;
23424: waveform_sig_loopback =-6415;
23425: waveform_sig_loopback =-8367;
23426: waveform_sig_loopback =-6675;
23427: waveform_sig_loopback =-6417;
23428: waveform_sig_loopback =-8254;
23429: waveform_sig_loopback =-6637;
23430: waveform_sig_loopback =-7262;
23431: waveform_sig_loopback =-7154;
23432: waveform_sig_loopback =-7587;
23433: waveform_sig_loopback =-6256;
23434: waveform_sig_loopback =-7718;
23435: waveform_sig_loopback =-7532;
23436: waveform_sig_loopback =-6467;
23437: waveform_sig_loopback =-7082;
23438: waveform_sig_loopback =-7924;
23439: waveform_sig_loopback =-6891;
23440: waveform_sig_loopback =-5913;
23441: waveform_sig_loopback =-8768;
23442: waveform_sig_loopback =-6886;
23443: waveform_sig_loopback =-5715;
23444: waveform_sig_loopback =-8248;
23445: waveform_sig_loopback =-7556;
23446: waveform_sig_loopback =-6006;
23447: waveform_sig_loopback =-6864;
23448: waveform_sig_loopback =-8296;
23449: waveform_sig_loopback =-6772;
23450: waveform_sig_loopback =-5766;
23451: waveform_sig_loopback =-8599;
23452: waveform_sig_loopback =-5052;
23453: waveform_sig_loopback =-8776;
23454: waveform_sig_loopback =-8574;
23455: waveform_sig_loopback =-4254;
23456: waveform_sig_loopback =-7072;
23457: waveform_sig_loopback =-7750;
23458: waveform_sig_loopback =-7987;
23459: waveform_sig_loopback =-6150;
23460: waveform_sig_loopback =-5552;
23461: waveform_sig_loopback =-7780;
23462: waveform_sig_loopback =-7531;
23463: waveform_sig_loopback =-6285;
23464: waveform_sig_loopback =-7121;
23465: waveform_sig_loopback =-6220;
23466: waveform_sig_loopback =-7998;
23467: waveform_sig_loopback =-6178;
23468: waveform_sig_loopback =-6308;
23469: waveform_sig_loopback =-7706;
23470: waveform_sig_loopback =-6099;
23471: waveform_sig_loopback =-7174;
23472: waveform_sig_loopback =-6433;
23473: waveform_sig_loopback =-7268;
23474: waveform_sig_loopback =-5897;
23475: waveform_sig_loopback =-6977;
23476: waveform_sig_loopback =-7474;
23477: waveform_sig_loopback =-5635;
23478: waveform_sig_loopback =-6721;
23479: waveform_sig_loopback =-7635;
23480: waveform_sig_loopback =-5766;
23481: waveform_sig_loopback =-6045;
23482: waveform_sig_loopback =-7979;
23483: waveform_sig_loopback =-5990;
23484: waveform_sig_loopback =-5562;
23485: waveform_sig_loopback =-7537;
23486: waveform_sig_loopback =-7009;
23487: waveform_sig_loopback =-5290;
23488: waveform_sig_loopback =-6204;
23489: waveform_sig_loopback =-7868;
23490: waveform_sig_loopback =-5948;
23491: waveform_sig_loopback =-5033;
23492: waveform_sig_loopback =-7849;
23493: waveform_sig_loopback =-4435;
23494: waveform_sig_loopback =-8249;
23495: waveform_sig_loopback =-7761;
23496: waveform_sig_loopback =-3193;
23497: waveform_sig_loopback =-6586;
23498: waveform_sig_loopback =-7389;
23499: waveform_sig_loopback =-6785;
23500: waveform_sig_loopback =-5536;
23501: waveform_sig_loopback =-4782;
23502: waveform_sig_loopback =-7058;
23503: waveform_sig_loopback =-6865;
23504: waveform_sig_loopback =-5147;
23505: waveform_sig_loopback =-6397;
23506: waveform_sig_loopback =-5548;
23507: waveform_sig_loopback =-6883;
23508: waveform_sig_loopback =-5410;
23509: waveform_sig_loopback =-5588;
23510: waveform_sig_loopback =-6621;
23511: waveform_sig_loopback =-5529;
23512: waveform_sig_loopback =-6034;
23513: waveform_sig_loopback =-5541;
23514: waveform_sig_loopback =-6683;
23515: waveform_sig_loopback =-4489;
23516: waveform_sig_loopback =-6362;
23517: waveform_sig_loopback =-6456;
23518: waveform_sig_loopback =-4389;
23519: waveform_sig_loopback =-6168;
23520: waveform_sig_loopback =-6325;
23521: waveform_sig_loopback =-4738;
23522: waveform_sig_loopback =-5396;
23523: waveform_sig_loopback =-6584;
23524: waveform_sig_loopback =-5101;
23525: waveform_sig_loopback =-4623;
23526: waveform_sig_loopback =-6261;
23527: waveform_sig_loopback =-6202;
23528: waveform_sig_loopback =-4026;
23529: waveform_sig_loopback =-5174;
23530: waveform_sig_loopback =-7038;
23531: waveform_sig_loopback =-4458;
23532: waveform_sig_loopback =-4139;
23533: waveform_sig_loopback =-6823;
23534: waveform_sig_loopback =-2956;
23535: waveform_sig_loopback =-7547;
23536: waveform_sig_loopback =-6348;
23537: waveform_sig_loopback =-1883;
23538: waveform_sig_loopback =-5860;
23539: waveform_sig_loopback =-5934;
23540: waveform_sig_loopback =-5585;
23541: waveform_sig_loopback =-4577;
23542: waveform_sig_loopback =-3190;
23543: waveform_sig_loopback =-6201;
23544: waveform_sig_loopback =-5537;
23545: waveform_sig_loopback =-3697;
23546: waveform_sig_loopback =-5566;
23547: waveform_sig_loopback =-3986;
23548: waveform_sig_loopback =-5705;
23549: waveform_sig_loopback =-4326;
23550: waveform_sig_loopback =-4033;
23551: waveform_sig_loopback =-5527;
23552: waveform_sig_loopback =-4252;
23553: waveform_sig_loopback =-4519;
23554: waveform_sig_loopback =-4524;
23555: waveform_sig_loopback =-5154;
23556: waveform_sig_loopback =-3096;
23557: waveform_sig_loopback =-5398;
23558: waveform_sig_loopback =-4730;
23559: waveform_sig_loopback =-3170;
23560: waveform_sig_loopback =-5029;
23561: waveform_sig_loopback =-4613;
23562: waveform_sig_loopback =-3587;
23563: waveform_sig_loopback =-3989;
23564: waveform_sig_loopback =-4989;
23565: waveform_sig_loopback =-3985;
23566: waveform_sig_loopback =-2986;
23567: waveform_sig_loopback =-4960;
23568: waveform_sig_loopback =-4878;
23569: waveform_sig_loopback =-2220;
23570: waveform_sig_loopback =-4082;
23571: waveform_sig_loopback =-5538;
23572: waveform_sig_loopback =-2613;
23573: waveform_sig_loopback =-3207;
23574: waveform_sig_loopback =-4985;
23575: waveform_sig_loopback =-1493;
23576: waveform_sig_loopback =-6561;
23577: waveform_sig_loopback =-4178;
23578: waveform_sig_loopback =-732;
23579: waveform_sig_loopback =-4397;
23580: waveform_sig_loopback =-4141;
23581: waveform_sig_loopback =-4442;
23582: waveform_sig_loopback =-2695;
23583: waveform_sig_loopback =-1676;
23584: waveform_sig_loopback =-5053;
23585: waveform_sig_loopback =-3488;
23586: waveform_sig_loopback =-2429;
23587: waveform_sig_loopback =-3974;
23588: waveform_sig_loopback =-2208;
23589: waveform_sig_loopback =-4449;
23590: waveform_sig_loopback =-2443;
23591: waveform_sig_loopback =-2480;
23592: waveform_sig_loopback =-4123;
23593: waveform_sig_loopback =-2439;
23594: waveform_sig_loopback =-2909;
23595: waveform_sig_loopback =-3160;
23596: waveform_sig_loopback =-3196;
23597: waveform_sig_loopback =-1664;
23598: waveform_sig_loopback =-3923;
23599: waveform_sig_loopback =-2574;
23600: waveform_sig_loopback =-2031;
23601: waveform_sig_loopback =-3085;
23602: waveform_sig_loopback =-2928;
23603: waveform_sig_loopback =-2193;
23604: waveform_sig_loopback =-1903;
23605: waveform_sig_loopback =-3754;
23606: waveform_sig_loopback =-2061;
23607: waveform_sig_loopback =-1111;
23608: waveform_sig_loopback =-3703;
23609: waveform_sig_loopback =-2793;
23610: waveform_sig_loopback =-619;
23611: waveform_sig_loopback =-2590;
23612: waveform_sig_loopback =-3569;
23613: waveform_sig_loopback =-947;
23614: waveform_sig_loopback =-1663;
23615: waveform_sig_loopback =-2988;
23616: waveform_sig_loopback =89;
23617: waveform_sig_loopback =-5009;
23618: waveform_sig_loopback =-1934;
23619: waveform_sig_loopback =642;
23620: waveform_sig_loopback =-2473;
23621: waveform_sig_loopback =-2386;
23622: waveform_sig_loopback =-2965;
23623: waveform_sig_loopback =-376;
23624: waveform_sig_loopback =-311;
23625: waveform_sig_loopback =-3344;
23626: waveform_sig_loopback =-1343;
23627: waveform_sig_loopback =-1130;
23628: waveform_sig_loopback =-1804;
23629: waveform_sig_loopback =-523;
23630: waveform_sig_loopback =-2944;
23631: waveform_sig_loopback =-140;
23632: waveform_sig_loopback =-1097;
23633: waveform_sig_loopback =-2239;
23634: waveform_sig_loopback =-373;
23635: waveform_sig_loopback =-1426;
23636: waveform_sig_loopback =-1134;
23637: waveform_sig_loopback =-1307;
23638: waveform_sig_loopback =-84;
23639: waveform_sig_loopback =-1827;
23640: waveform_sig_loopback =-897;
23641: waveform_sig_loopback =-280;
23642: waveform_sig_loopback =-1004;
23643: waveform_sig_loopback =-1368;
23644: waveform_sig_loopback =-156;
23645: waveform_sig_loopback =-21;
23646: waveform_sig_loopback =-2188;
23647: waveform_sig_loopback =138;
23648: waveform_sig_loopback =542;
23649: waveform_sig_loopback =-2040;
23650: waveform_sig_loopback =-547;
23651: waveform_sig_loopback =995;
23652: waveform_sig_loopback =-764;
23653: waveform_sig_loopback =-1487;
23654: waveform_sig_loopback =731;
23655: waveform_sig_loopback =301;
23656: waveform_sig_loopback =-1023;
23657: waveform_sig_loopback =1700;
23658: waveform_sig_loopback =-2958;
23659: waveform_sig_loopback =-8;
23660: waveform_sig_loopback =2363;
23661: waveform_sig_loopback =-388;
23662: waveform_sig_loopback =-847;
23663: waveform_sig_loopback =-781;
23664: waveform_sig_loopback =1602;
23665: waveform_sig_loopback =1154;
23666: waveform_sig_loopback =-1086;
23667: waveform_sig_loopback =417;
23668: waveform_sig_loopback =637;
23669: waveform_sig_loopback =443;
23670: waveform_sig_loopback =931;
23671: waveform_sig_loopback =-756;
23672: waveform_sig_loopback =1843;
23673: waveform_sig_loopback =428;
23674: waveform_sig_loopback =80;
23675: waveform_sig_loopback =1274;
23676: waveform_sig_loopback =433;
23677: waveform_sig_loopback =940;
23678: waveform_sig_loopback =378;
23679: waveform_sig_loopback =1929;
23680: waveform_sig_loopback =59;
23681: waveform_sig_loopback =829;
23682: waveform_sig_loopback =1825;
23683: waveform_sig_loopback =776;
23684: waveform_sig_loopback =393;
23685: waveform_sig_loopback =2021;
23686: waveform_sig_loopback =1576;
23687: waveform_sig_loopback =-307;
23688: waveform_sig_loopback =2320;
23689: waveform_sig_loopback =2095;
23690: waveform_sig_loopback =-59;
23691: waveform_sig_loopback =1559;
23692: waveform_sig_loopback =2516;
23693: waveform_sig_loopback =1375;
23694: waveform_sig_loopback =230;
23695: waveform_sig_loopback =2550;
23696: waveform_sig_loopback =2444;
23697: waveform_sig_loopback =527;
23698: waveform_sig_loopback =3748;
23699: waveform_sig_loopback =-1177;
23700: waveform_sig_loopback =1790;
23701: waveform_sig_loopback =4557;
23702: waveform_sig_loopback =1063;
23703: waveform_sig_loopback =934;
23704: waveform_sig_loopback =1506;
23705: waveform_sig_loopback =3099;
23706: waveform_sig_loopback =3141;
23707: waveform_sig_loopback =791;
23708: waveform_sig_loopback =2103;
23709: waveform_sig_loopback =2749;
23710: waveform_sig_loopback =2138;
23711: waveform_sig_loopback =2645;
23712: waveform_sig_loopback =1374;
23713: waveform_sig_loopback =3465;
23714: waveform_sig_loopback =2231;
23715: waveform_sig_loopback =2082;
23716: waveform_sig_loopback =2929;
23717: waveform_sig_loopback =2457;
23718: waveform_sig_loopback =2737;
23719: waveform_sig_loopback =2058;
23720: waveform_sig_loopback =3988;
23721: waveform_sig_loopback =1746;
23722: waveform_sig_loopback =2582;
23723: waveform_sig_loopback =3938;
23724: waveform_sig_loopback =2207;
23725: waveform_sig_loopback =2379;
23726: waveform_sig_loopback =4110;
23727: waveform_sig_loopback =2804;
23728: waveform_sig_loopback =2024;
23729: waveform_sig_loopback =3988;
23730: waveform_sig_loopback =3634;
23731: waveform_sig_loopback =2084;
23732: waveform_sig_loopback =3001;
23733: waveform_sig_loopback =4596;
23734: waveform_sig_loopback =3053;
23735: waveform_sig_loopback =1741;
23736: waveform_sig_loopback =4858;
23737: waveform_sig_loopback =3790;
23738: waveform_sig_loopback =2347;
23739: waveform_sig_loopback =5721;
23740: waveform_sig_loopback =138;
23741: waveform_sig_loopback =3996;
23742: waveform_sig_loopback =6192;
23743: waveform_sig_loopback =2579;
23744: waveform_sig_loopback =2934;
23745: waveform_sig_loopback =3232;
23746: waveform_sig_loopback =4787;
23747: waveform_sig_loopback =4927;
23748: waveform_sig_loopback =2334;
23749: waveform_sig_loopback =3948;
23750: waveform_sig_loopback =4543;
23751: waveform_sig_loopback =3656;
23752: waveform_sig_loopback =4322;
23753: waveform_sig_loopback =3266;
23754: waveform_sig_loopback =4882;
23755: waveform_sig_loopback =4125;
23756: waveform_sig_loopback =3752;
23757: waveform_sig_loopback =4272;
23758: waveform_sig_loopback =4607;
23759: waveform_sig_loopback =3882;
23760: waveform_sig_loopback =3963;
23761: waveform_sig_loopback =5816;
23762: waveform_sig_loopback =2814;
23763: waveform_sig_loopback =4876;
23764: waveform_sig_loopback =5206;
23765: waveform_sig_loopback =3784;
23766: waveform_sig_loopback =4351;
23767: waveform_sig_loopback =5320;
23768: waveform_sig_loopback =4604;
23769: waveform_sig_loopback =3617;
23770: waveform_sig_loopback =5458;
23771: waveform_sig_loopback =5393;
23772: waveform_sig_loopback =3523;
23773: waveform_sig_loopback =4584;
23774: waveform_sig_loopback =6367;
23775: waveform_sig_loopback =4377;
23776: waveform_sig_loopback =3330;
23777: waveform_sig_loopback =6733;
23778: waveform_sig_loopback =4883;
23779: waveform_sig_loopback =4216;
23780: waveform_sig_loopback =7233;
23781: waveform_sig_loopback =1256;
23782: waveform_sig_loopback =6101;
23783: waveform_sig_loopback =7432;
23784: waveform_sig_loopback =3903;
23785: waveform_sig_loopback =4704;
23786: waveform_sig_loopback =4396;
23787: waveform_sig_loopback =6451;
23788: waveform_sig_loopback =6507;
23789: waveform_sig_loopback =3400;
23790: waveform_sig_loopback =5778;
23791: waveform_sig_loopback =5826;
23792: waveform_sig_loopback =4941;
23793: waveform_sig_loopback =6141;
23794: waveform_sig_loopback =4228;
23795: waveform_sig_loopback =6463;
23796: waveform_sig_loopback =5658;
23797: waveform_sig_loopback =4750;
23798: waveform_sig_loopback =5988;
23799: waveform_sig_loopback =5639;
23800: waveform_sig_loopback =5198;
23801: waveform_sig_loopback =5840;
23802: waveform_sig_loopback =6512;
23803: waveform_sig_loopback =4148;
23804: waveform_sig_loopback =6534;
23805: waveform_sig_loopback =6236;
23806: waveform_sig_loopback =5250;
23807: waveform_sig_loopback =5358;
23808: waveform_sig_loopback =6703;
23809: waveform_sig_loopback =6074;
23810: waveform_sig_loopback =4582;
23811: waveform_sig_loopback =6830;
23812: waveform_sig_loopback =6626;
23813: waveform_sig_loopback =4690;
23814: waveform_sig_loopback =5818;
23815: waveform_sig_loopback =7590;
23816: waveform_sig_loopback =5366;
23817: waveform_sig_loopback =4693;
23818: waveform_sig_loopback =7990;
23819: waveform_sig_loopback =5508;
23820: waveform_sig_loopback =6035;
23821: waveform_sig_loopback =7970;
23822: waveform_sig_loopback =2170;
23823: waveform_sig_loopback =7882;
23824: waveform_sig_loopback =7897;
23825: waveform_sig_loopback =5376;
23826: waveform_sig_loopback =5687;
23827: waveform_sig_loopback =5203;
23828: waveform_sig_loopback =8191;
23829: waveform_sig_loopback =6996;
23830: waveform_sig_loopback =4503;
23831: waveform_sig_loopback =7247;
23832: waveform_sig_loopback =6322;
23833: waveform_sig_loopback =6482;
23834: waveform_sig_loopback =6898;
23835: waveform_sig_loopback =5121;
23836: waveform_sig_loopback =8040;
23837: waveform_sig_loopback =6073;
23838: waveform_sig_loopback =5980;
23839: waveform_sig_loopback =7161;
23840: waveform_sig_loopback =6511;
23841: waveform_sig_loopback =6251;
23842: waveform_sig_loopback =6655;
23843: waveform_sig_loopback =7528;
23844: waveform_sig_loopback =5376;
23845: waveform_sig_loopback =7284;
23846: waveform_sig_loopback =6949;
23847: waveform_sig_loopback =6374;
23848: waveform_sig_loopback =6412;
23849: waveform_sig_loopback =7382;
23850: waveform_sig_loopback =6985;
23851: waveform_sig_loopback =5391;
23852: waveform_sig_loopback =7893;
23853: waveform_sig_loopback =7498;
23854: waveform_sig_loopback =5057;
23855: waveform_sig_loopback =7288;
23856: waveform_sig_loopback =8197;
23857: waveform_sig_loopback =5846;
23858: waveform_sig_loopback =6035;
23859: waveform_sig_loopback =8337;
23860: waveform_sig_loopback =6567;
23861: waveform_sig_loopback =6852;
23862: waveform_sig_loopback =8188;
23863: waveform_sig_loopback =3599;
23864: waveform_sig_loopback =8327;
23865: waveform_sig_loopback =8515;
23866: waveform_sig_loopback =6442;
23867: waveform_sig_loopback =5893;
23868: waveform_sig_loopback =6360;
23869: waveform_sig_loopback =8733;
23870: waveform_sig_loopback =7412;
23871: waveform_sig_loopback =5591;
23872: waveform_sig_loopback =7588;
23873: waveform_sig_loopback =6954;
23874: waveform_sig_loopback =7320;
23875: waveform_sig_loopback =7211;
23876: waveform_sig_loopback =5886;
23877: waveform_sig_loopback =8625;
23878: waveform_sig_loopback =6446;
23879: waveform_sig_loopback =6840;
23880: waveform_sig_loopback =7583;
23881: waveform_sig_loopback =6915;
23882: waveform_sig_loopback =6998;
23883: waveform_sig_loopback =7115;
23884: waveform_sig_loopback =7923;
23885: waveform_sig_loopback =6021;
23886: waveform_sig_loopback =7572;
23887: waveform_sig_loopback =7543;
23888: waveform_sig_loopback =6904;
23889: waveform_sig_loopback =6505;
23890: waveform_sig_loopback =8275;
23891: waveform_sig_loopback =7137;
23892: waveform_sig_loopback =5717;
23893: waveform_sig_loopback =8741;
23894: waveform_sig_loopback =7336;
23895: waveform_sig_loopback =5715;
23896: waveform_sig_loopback =7828;
23897: waveform_sig_loopback =8119;
23898: waveform_sig_loopback =6622;
23899: waveform_sig_loopback =6121;
23900: waveform_sig_loopback =8682;
23901: waveform_sig_loopback =7119;
23902: waveform_sig_loopback =6851;
23903: waveform_sig_loopback =8636;
23904: waveform_sig_loopback =3820;
23905: waveform_sig_loopback =8547;
23906: waveform_sig_loopback =9064;
23907: waveform_sig_loopback =6277;
23908: waveform_sig_loopback =6145;
23909: waveform_sig_loopback =6958;
23910: waveform_sig_loopback =8555;
23911: waveform_sig_loopback =7773;
23912: waveform_sig_loopback =5723;
23913: waveform_sig_loopback =7679;
23914: waveform_sig_loopback =7276;
23915: waveform_sig_loopback =7348;
23916: waveform_sig_loopback =7258;
23917: waveform_sig_loopback =6270;
23918: waveform_sig_loopback =8591;
23919: waveform_sig_loopback =6437;
23920: waveform_sig_loopback =7135;
23921: waveform_sig_loopback =7478;
23922: waveform_sig_loopback =7001;
23923: waveform_sig_loopback =7115;
23924: waveform_sig_loopback =6960;
23925: waveform_sig_loopback =8127;
23926: waveform_sig_loopback =6006;
23927: waveform_sig_loopback =7303;
23928: waveform_sig_loopback =8026;
23929: waveform_sig_loopback =6334;
23930: waveform_sig_loopback =6755;
23931: waveform_sig_loopback =8423;
23932: waveform_sig_loopback =6386;
23933: waveform_sig_loopback =6326;
23934: waveform_sig_loopback =8303;
23935: waveform_sig_loopback =7165;
23936: waveform_sig_loopback =5956;
23937: waveform_sig_loopback =7329;
23938: waveform_sig_loopback =8288;
23939: waveform_sig_loopback =6283;
23940: waveform_sig_loopback =5874;
23941: waveform_sig_loopback =8827;
23942: waveform_sig_loopback =6522;
23943: waveform_sig_loopback =6786;
23944: waveform_sig_loopback =8434;
23945: waveform_sig_loopback =3384;
23946: waveform_sig_loopback =8567;
23947: waveform_sig_loopback =8758;
23948: waveform_sig_loopback =5835;
23949: waveform_sig_loopback =6037;
23950: waveform_sig_loopback =6706;
23951: waveform_sig_loopback =8150;
23952: waveform_sig_loopback =7572;
23953: waveform_sig_loopback =5299;
23954: waveform_sig_loopback =7311;
23955: waveform_sig_loopback =7149;
23956: waveform_sig_loopback =6803;
23957: waveform_sig_loopback =6928;
23958: waveform_sig_loopback =6070;
23959: waveform_sig_loopback =7942;
23960: waveform_sig_loopback =6255;
23961: waveform_sig_loopback =6683;
23962: waveform_sig_loopback =6842;
23963: waveform_sig_loopback =6989;
23964: waveform_sig_loopback =6285;
23965: waveform_sig_loopback =6686;
23966: waveform_sig_loopback =7798;
23967: waveform_sig_loopback =5113;
23968: waveform_sig_loopback =7324;
23969: waveform_sig_loopback =7299;
23970: waveform_sig_loopback =5700;
23971: waveform_sig_loopback =6640;
23972: waveform_sig_loopback =7540;
23973: waveform_sig_loopback =5955;
23974: waveform_sig_loopback =5936;
23975: waveform_sig_loopback =7486;
23976: waveform_sig_loopback =6769;
23977: waveform_sig_loopback =5289;
23978: waveform_sig_loopback =6647;
23979: waveform_sig_loopback =7912;
23980: waveform_sig_loopback =5392;
23981: waveform_sig_loopback =5347;
23982: waveform_sig_loopback =8410;
23983: waveform_sig_loopback =5446;
23984: waveform_sig_loopback =6592;
23985: waveform_sig_loopback =7545;
23986: waveform_sig_loopback =2480;
23987: waveform_sig_loopback =8426;
23988: waveform_sig_loopback =7692;
23989: waveform_sig_loopback =5060;
23990: waveform_sig_loopback =5516;
23991: waveform_sig_loopback =5734;
23992: waveform_sig_loopback =7624;
23993: waveform_sig_loopback =6763;
23994: waveform_sig_loopback =4220;
23995: waveform_sig_loopback =6909;
23996: waveform_sig_loopback =6128;
23997: waveform_sig_loopback =5958;
23998: waveform_sig_loopback =6244;
23999: waveform_sig_loopback =5022;
24000: waveform_sig_loopback =7211;
24001: waveform_sig_loopback =5462;
24002: waveform_sig_loopback =5595;
24003: waveform_sig_loopback =6124;
24004: waveform_sig_loopback =6093;
24005: waveform_sig_loopback =5084;
24006: waveform_sig_loopback =6206;
24007: waveform_sig_loopback =6555;
24008: waveform_sig_loopback =4137;
24009: waveform_sig_loopback =6769;
24010: waveform_sig_loopback =5842;
24011: waveform_sig_loopback =4984;
24012: waveform_sig_loopback =5708;
24013: waveform_sig_loopback =6248;
24014: waveform_sig_loopback =5329;
24015: waveform_sig_loopback =4662;
24016: waveform_sig_loopback =6511;
24017: waveform_sig_loopback =5901;
24018: waveform_sig_loopback =3855;
24019: waveform_sig_loopback =5952;
24020: waveform_sig_loopback =6790;
24021: waveform_sig_loopback =4021;
24022: waveform_sig_loopback =4677;
24023: waveform_sig_loopback =7128;
24024: waveform_sig_loopback =4220;
24025: waveform_sig_loopback =5866;
24026: waveform_sig_loopback =5974;
24027: waveform_sig_loopback =1518;
24028: waveform_sig_loopback =7564;
24029: waveform_sig_loopback =6179;
24030: waveform_sig_loopback =4087;
24031: waveform_sig_loopback =4336;
24032: waveform_sig_loopback =4421;
24033: waveform_sig_loopback =6779;
24034: waveform_sig_loopback =5274;
24035: waveform_sig_loopback =2997;
24036: waveform_sig_loopback =6052;
24037: waveform_sig_loopback =4452;
24038: waveform_sig_loopback =5038;
24039: waveform_sig_loopback =4949;
24040: waveform_sig_loopback =3519;
24041: waveform_sig_loopback =6344;
24042: waveform_sig_loopback =3859;
24043: waveform_sig_loopback =4329;
24044: waveform_sig_loopback =5109;
24045: waveform_sig_loopback =4426;
24046: waveform_sig_loopback =3978;
24047: waveform_sig_loopback =5036;
24048: waveform_sig_loopback =4778;
24049: waveform_sig_loopback =3226;
24050: waveform_sig_loopback =5243;
24051: waveform_sig_loopback =4341;
24052: waveform_sig_loopback =3930;
24053: waveform_sig_loopback =4044;
24054: waveform_sig_loopback =5052;
24055: waveform_sig_loopback =3924;
24056: waveform_sig_loopback =3027;
24057: waveform_sig_loopback =5500;
24058: waveform_sig_loopback =4217;
24059: waveform_sig_loopback =2317;
24060: waveform_sig_loopback =4957;
24061: waveform_sig_loopback =4957;
24062: waveform_sig_loopback =2671;
24063: waveform_sig_loopback =3391;
24064: waveform_sig_loopback =5452;
24065: waveform_sig_loopback =2881;
24066: waveform_sig_loopback =4447;
24067: waveform_sig_loopback =4215;
24068: waveform_sig_loopback =240;
24069: waveform_sig_loopback =6160;
24070: waveform_sig_loopback =4447;
24071: waveform_sig_loopback =2727;
24072: waveform_sig_loopback =2630;
24073: waveform_sig_loopback =3009;
24074: waveform_sig_loopback =5445;
24075: waveform_sig_loopback =3261;
24076: waveform_sig_loopback =1782;
24077: waveform_sig_loopback =4508;
24078: waveform_sig_loopback =2553;
24079: waveform_sig_loopback =3963;
24080: waveform_sig_loopback =2897;
24081: waveform_sig_loopback =2191;
24082: waveform_sig_loopback =4942;
24083: waveform_sig_loopback =1753;
24084: waveform_sig_loopback =3255;
24085: waveform_sig_loopback =3297;
24086: waveform_sig_loopback =2651;
24087: waveform_sig_loopback =2765;
24088: waveform_sig_loopback =3017;
24089: waveform_sig_loopback =3339;
24090: waveform_sig_loopback =1701;
24091: waveform_sig_loopback =3263;
24092: waveform_sig_loopback =3095;
24093: waveform_sig_loopback =1974;
24094: waveform_sig_loopback =2470;
24095: waveform_sig_loopback =3627;
24096: waveform_sig_loopback =1839;
24097: waveform_sig_loopback =1643;
24098: waveform_sig_loopback =3831;
24099: waveform_sig_loopback =2422;
24100: waveform_sig_loopback =701;
24101: waveform_sig_loopback =3398;
24102: waveform_sig_loopback =3069;
24103: waveform_sig_loopback =1026;
24104: waveform_sig_loopback =1818;
24105: waveform_sig_loopback =3508;
24106: waveform_sig_loopback =1365;
24107: waveform_sig_loopback =2717;
24108: waveform_sig_loopback =2156;
24109: waveform_sig_loopback =-1078;
24110: waveform_sig_loopback =4160;
24111: waveform_sig_loopback =2770;
24112: waveform_sig_loopback =1092;
24113: waveform_sig_loopback =467;
24114: waveform_sig_loopback =1862;
24115: waveform_sig_loopback =3352;
24116: waveform_sig_loopback =1347;
24117: waveform_sig_loopback =498;
24118: waveform_sig_loopback =2153;
24119: waveform_sig_loopback =1280;
24120: waveform_sig_loopback =2113;
24121: waveform_sig_loopback =719;
24122: waveform_sig_loopback =1106;
24123: waveform_sig_loopback =2551;
24124: waveform_sig_loopback =177;
24125: waveform_sig_loopback =1640;
24126: waveform_sig_loopback =1048;
24127: waveform_sig_loopback =1317;
24128: waveform_sig_loopback =632;
24129: waveform_sig_loopback =1382;
24130: waveform_sig_loopback =1518;
24131: waveform_sig_loopback =-247;
24132: waveform_sig_loopback =1653;
24133: waveform_sig_loopback =1138;
24134: waveform_sig_loopback =126;
24135: waveform_sig_loopback =559;
24136: waveform_sig_loopback =1935;
24137: waveform_sig_loopback =-254;
24138: waveform_sig_loopback =-74;
24139: waveform_sig_loopback =2131;
24140: waveform_sig_loopback =25;
24141: waveform_sig_loopback =-648;
24142: waveform_sig_loopback =1357;
24143: waveform_sig_loopback =1058;
24144: waveform_sig_loopback =-547;
24145: waveform_sig_loopback =-405;
24146: waveform_sig_loopback =2011;
24147: waveform_sig_loopback =-617;
24148: waveform_sig_loopback =713;
24149: waveform_sig_loopback =537;
24150: waveform_sig_loopback =-3346;
24151: waveform_sig_loopback =2621;
24152: waveform_sig_loopback =1146;
24153: waveform_sig_loopback =-1379;
24154: waveform_sig_loopback =-1143;
24155: waveform_sig_loopback =33;
24156: waveform_sig_loopback =1338;
24157: waveform_sig_loopback =-207;
24158: waveform_sig_loopback =-1850;
24159: waveform_sig_loopback =429;
24160: waveform_sig_loopback =-321;
24161: waveform_sig_loopback =-233;
24162: waveform_sig_loopback =-954;
24163: waveform_sig_loopback =-832;
24164: waveform_sig_loopback =498;
24165: waveform_sig_loopback =-1490;
24166: waveform_sig_loopback =-618;
24167: waveform_sig_loopback =-678;
24168: waveform_sig_loopback =-517;
24169: waveform_sig_loopback =-1525;
24170: waveform_sig_loopback =-420;
24171: waveform_sig_loopback =-445;
24172: waveform_sig_loopback =-2160;
24173: waveform_sig_loopback =-279;
24174: waveform_sig_loopback =-700;
24175: waveform_sig_loopback =-1956;
24176: waveform_sig_loopback =-1000;
24177: waveform_sig_loopback =-94;
24178: waveform_sig_loopback =-2437;
24179: waveform_sig_loopback =-1377;
24180: waveform_sig_loopback =-138;
24181: waveform_sig_loopback =-1810;
24182: waveform_sig_loopback =-2301;
24183: waveform_sig_loopback =-876;
24184: waveform_sig_loopback =-341;
24185: waveform_sig_loopback =-2855;
24186: waveform_sig_loopback =-2240;
24187: waveform_sig_loopback =606;
24188: waveform_sig_loopback =-3287;
24189: waveform_sig_loopback =-561;
24190: waveform_sig_loopback =-1688;
24191: waveform_sig_loopback =-5242;
24192: waveform_sig_loopback =1252;
24193: waveform_sig_loopback =-1526;
24194: waveform_sig_loopback =-3050;
24195: waveform_sig_loopback =-2634;
24196: waveform_sig_loopback =-2238;
24197: waveform_sig_loopback =-412;
24198: waveform_sig_loopback =-2339;
24199: waveform_sig_loopback =-3633;
24200: waveform_sig_loopback =-1201;
24201: waveform_sig_loopback =-2674;
24202: waveform_sig_loopback =-1980;
24203: waveform_sig_loopback =-2699;
24204: waveform_sig_loopback =-2763;
24205: waveform_sig_loopback =-1428;
24206: waveform_sig_loopback =-3284;
24207: waveform_sig_loopback =-2415;
24208: waveform_sig_loopback =-2582;
24209: waveform_sig_loopback =-2256;
24210: waveform_sig_loopback =-3595;
24211: waveform_sig_loopback =-1852;
24212: waveform_sig_loopback =-2474;
24213: waveform_sig_loopback =-4210;
24214: waveform_sig_loopback =-1468;
24215: waveform_sig_loopback =-3018;
24216: waveform_sig_loopback =-3577;
24217: waveform_sig_loopback =-2594;
24218: waveform_sig_loopback =-2431;
24219: waveform_sig_loopback =-3686;
24220: waveform_sig_loopback =-3536;
24221: waveform_sig_loopback =-1968;
24222: waveform_sig_loopback =-3308;
24223: waveform_sig_loopback =-4585;
24224: waveform_sig_loopback =-2258;
24225: waveform_sig_loopback =-2328;
24226: waveform_sig_loopback =-4907;
24227: waveform_sig_loopback =-3505;
24228: waveform_sig_loopback =-1579;
24229: waveform_sig_loopback =-5054;
24230: waveform_sig_loopback =-1964;
24231: waveform_sig_loopback =-4024;
24232: waveform_sig_loopback =-6650;
24233: waveform_sig_loopback =-421;
24234: waveform_sig_loopback =-3577;
24235: waveform_sig_loopback =-4541;
24236: waveform_sig_loopback =-4541;
24237: waveform_sig_loopback =-3933;
24238: waveform_sig_loopback =-1850;
24239: waveform_sig_loopback =-4355;
24240: waveform_sig_loopback =-5306;
24241: waveform_sig_loopback =-2714;
24242: waveform_sig_loopback =-4583;
24243: waveform_sig_loopback =-3440;
24244: waveform_sig_loopback =-4461;
24245: waveform_sig_loopback =-4562;
24246: waveform_sig_loopback =-2808;
24247: waveform_sig_loopback =-5107;
24248: waveform_sig_loopback =-4129;
24249: waveform_sig_loopback =-3962;
24250: waveform_sig_loopback =-4200;
24251: waveform_sig_loopback =-5127;
24252: waveform_sig_loopback =-3219;
24253: waveform_sig_loopback =-4623;
24254: waveform_sig_loopback =-5369;
24255: waveform_sig_loopback =-3292;
24256: waveform_sig_loopback =-4871;
24257: waveform_sig_loopback =-4788;
24258: waveform_sig_loopback =-4653;
24259: waveform_sig_loopback =-3717;
24260: waveform_sig_loopback =-5300;
24261: waveform_sig_loopback =-5367;
24262: waveform_sig_loopback =-3165;
24263: waveform_sig_loopback =-5224;
24264: waveform_sig_loopback =-6099;
24265: waveform_sig_loopback =-3565;
24266: waveform_sig_loopback =-4169;
24267: waveform_sig_loopback =-6404;
24268: waveform_sig_loopback =-4839;
24269: waveform_sig_loopback =-3349;
24270: waveform_sig_loopback =-6467;
24271: waveform_sig_loopback =-3339;
24272: waveform_sig_loopback =-5975;
24273: waveform_sig_loopback =-7693;
24274: waveform_sig_loopback =-1993;
24275: waveform_sig_loopback =-5208;
24276: waveform_sig_loopback =-5779;
24277: waveform_sig_loopback =-6300;
24278: waveform_sig_loopback =-5110;
24279: waveform_sig_loopback =-3262;
24280: waveform_sig_loopback =-6199;
24281: waveform_sig_loopback =-6330;
24282: waveform_sig_loopback =-4264;
24283: waveform_sig_loopback =-6148;
24284: waveform_sig_loopback =-4473;
24285: waveform_sig_loopback =-6290;
24286: waveform_sig_loopback =-5744;
24287: waveform_sig_loopback =-4080;
24288: waveform_sig_loopback =-6848;
24289: waveform_sig_loopback =-5142;
24290: waveform_sig_loopback =-5483;
24291: waveform_sig_loopback =-5721;
24292: waveform_sig_loopback =-6132;
24293: waveform_sig_loopback =-4932;
24294: waveform_sig_loopback =-5875;
24295: waveform_sig_loopback =-6501;
24296: waveform_sig_loopback =-5020;
24297: waveform_sig_loopback =-5821;
24298: waveform_sig_loopback =-6306;
24299: waveform_sig_loopback =-6027;
24300: waveform_sig_loopback =-4733;
24301: waveform_sig_loopback =-6979;
24302: waveform_sig_loopback =-6406;
24303: waveform_sig_loopback =-4396;
24304: waveform_sig_loopback =-6758;
24305: waveform_sig_loopback =-7074;
24306: waveform_sig_loopback =-4822;
24307: waveform_sig_loopback =-5647;
24308: waveform_sig_loopback =-7440;
24309: waveform_sig_loopback =-6015;
24310: waveform_sig_loopback =-4743;
24311: waveform_sig_loopback =-7439;
24312: waveform_sig_loopback =-4591;
24313: waveform_sig_loopback =-7353;
24314: waveform_sig_loopback =-8456;
24315: waveform_sig_loopback =-3480;
24316: waveform_sig_loopback =-6132;
24317: waveform_sig_loopback =-6968;
24318: waveform_sig_loopback =-7674;
24319: waveform_sig_loopback =-5694;
24320: waveform_sig_loopback =-4804;
24321: waveform_sig_loopback =-7209;
24322: waveform_sig_loopback =-7160;
24323: waveform_sig_loopback =-5762;
24324: waveform_sig_loopback =-6783;
24325: waveform_sig_loopback =-5692;
24326: waveform_sig_loopback =-7487;
24327: waveform_sig_loopback =-6366;
24328: waveform_sig_loopback =-5524;
24329: waveform_sig_loopback =-7689;
24330: waveform_sig_loopback =-6045;
24331: waveform_sig_loopback =-6743;
24332: waveform_sig_loopback =-6451;
24333: waveform_sig_loopback =-7167;
24334: waveform_sig_loopback =-5944;
24335: waveform_sig_loopback =-6743;
24336: waveform_sig_loopback =-7447;
24337: waveform_sig_loopback =-5999;
24338: waveform_sig_loopback =-6575;
24339: waveform_sig_loopback =-7427;
24340: waveform_sig_loopback =-6744;
24341: waveform_sig_loopback =-5503;
24342: waveform_sig_loopback =-8200;
24343: waveform_sig_loopback =-6788;
24344: waveform_sig_loopback =-5405;
24345: waveform_sig_loopback =-7836;
24346: waveform_sig_loopback =-7410;
24347: waveform_sig_loopback =-5979;
24348: waveform_sig_loopback =-6291;
24349: waveform_sig_loopback =-8140;
24350: waveform_sig_loopback =-6983;
24351: waveform_sig_loopback =-5203;
24352: waveform_sig_loopback =-8453;
24353: waveform_sig_loopback =-5240;
24354: waveform_sig_loopback =-8121;
24355: waveform_sig_loopback =-9220;
24356: waveform_sig_loopback =-4009;
24357: waveform_sig_loopback =-6901;
24358: waveform_sig_loopback =-7963;
24359: waveform_sig_loopback =-8041;
24360: waveform_sig_loopback =-6337;
24361: waveform_sig_loopback =-5696;
24362: waveform_sig_loopback =-7662;
24363: waveform_sig_loopback =-7928;
24364: waveform_sig_loopback =-6357;
24365: waveform_sig_loopback =-7267;
24366: waveform_sig_loopback =-6619;
24367: waveform_sig_loopback =-7867;
24368: waveform_sig_loopback =-6879;
24369: waveform_sig_loopback =-6387;
24370: waveform_sig_loopback =-7966;
24371: waveform_sig_loopback =-6732;
24372: waveform_sig_loopback =-7298;
24373: waveform_sig_loopback =-6795;
24374: waveform_sig_loopback =-7937;
24375: waveform_sig_loopback =-6283;
24376: waveform_sig_loopback =-7219;
24377: waveform_sig_loopback =-8185;
24378: waveform_sig_loopback =-6115;
24379: waveform_sig_loopback =-7166;
24380: waveform_sig_loopback =-8038;
24381: waveform_sig_loopback =-6765;
24382: waveform_sig_loopback =-6423;
24383: waveform_sig_loopback =-8359;
24384: waveform_sig_loopback =-7012;
24385: waveform_sig_loopback =-6182;
24386: waveform_sig_loopback =-7938;
24387: waveform_sig_loopback =-7943;
24388: waveform_sig_loopback =-6278;
24389: waveform_sig_loopback =-6578;
24390: waveform_sig_loopback =-8669;
24391: waveform_sig_loopback =-7078;
24392: waveform_sig_loopback =-5531;
24393: waveform_sig_loopback =-8931;
24394: waveform_sig_loopback =-5295;
24395: waveform_sig_loopback =-8583;
24396: waveform_sig_loopback =-9505;
24397: waveform_sig_loopback =-3921;
24398: waveform_sig_loopback =-7386;
24399: waveform_sig_loopback =-8277;
24400: waveform_sig_loopback =-7946;
24401: waveform_sig_loopback =-6839;
24402: waveform_sig_loopback =-5692;
24403: waveform_sig_loopback =-7915;
24404: waveform_sig_loopback =-8293;
24405: waveform_sig_loopback =-6152;
24406: waveform_sig_loopback =-7636;
24407: waveform_sig_loopback =-6760;
24408: waveform_sig_loopback =-7835;
24409: waveform_sig_loopback =-7192;
24410: waveform_sig_loopback =-6380;
24411: waveform_sig_loopback =-8028;
24412: waveform_sig_loopback =-7003;
24413: waveform_sig_loopback =-7129;
24414: waveform_sig_loopback =-6981;
24415: waveform_sig_loopback =-8066;
24416: waveform_sig_loopback =-6033;
24417: waveform_sig_loopback =-7511;
24418: waveform_sig_loopback =-8070;
24419: waveform_sig_loopback =-5945;
24420: waveform_sig_loopback =-7512;
24421: waveform_sig_loopback =-7733;
24422: waveform_sig_loopback =-6629;
24423: waveform_sig_loopback =-6684;
24424: waveform_sig_loopback =-8049;
24425: waveform_sig_loopback =-7138;
24426: waveform_sig_loopback =-5992;
24427: waveform_sig_loopback =-7714;
24428: waveform_sig_loopback =-8068;
24429: waveform_sig_loopback =-5821;
24430: waveform_sig_loopback =-6642;
24431: waveform_sig_loopback =-8707;
24432: waveform_sig_loopback =-6593;
24433: waveform_sig_loopback =-5590;
24434: waveform_sig_loopback =-8736;
24435: waveform_sig_loopback =-4879;
24436: waveform_sig_loopback =-8794;
24437: waveform_sig_loopback =-8980;
24438: waveform_sig_loopback =-3600;
24439: waveform_sig_loopback =-7524;
24440: waveform_sig_loopback =-7791;
24441: waveform_sig_loopback =-7704;
24442: waveform_sig_loopback =-6697;
24443: waveform_sig_loopback =-5021;
24444: waveform_sig_loopback =-8018;
24445: waveform_sig_loopback =-7765;
24446: waveform_sig_loopback =-5728;
24447: waveform_sig_loopback =-7664;
24448: waveform_sig_loopback =-5983;
24449: waveform_sig_loopback =-7705;
24450: waveform_sig_loopback =-6784;
24451: waveform_sig_loopback =-5780;
24452: waveform_sig_loopback =-7893;
24453: waveform_sig_loopback =-6379;
24454: waveform_sig_loopback =-6698;
24455: waveform_sig_loopback =-6726;
24456: waveform_sig_loopback =-7403;
24457: waveform_sig_loopback =-5528;
24458: waveform_sig_loopback =-7257;
24459: waveform_sig_loopback =-7328;
24460: waveform_sig_loopback =-5534;
24461: waveform_sig_loopback =-7129;
24462: waveform_sig_loopback =-7017;
24463: waveform_sig_loopback =-6165;
24464: waveform_sig_loopback =-6115;
24465: waveform_sig_loopback =-7323;
24466: waveform_sig_loopback =-6689;
24467: waveform_sig_loopback =-5253;
24468: waveform_sig_loopback =-7177;
24469: waveform_sig_loopback =-7613;
24470: waveform_sig_loopback =-4819;
24471: waveform_sig_loopback =-6337;
24472: waveform_sig_loopback =-7963;
24473: waveform_sig_loopback =-5521;
24474: waveform_sig_loopback =-5508;
24475: waveform_sig_loopback =-7624;
24476: waveform_sig_loopback =-4193;
24477: waveform_sig_loopback =-8560;
24478: waveform_sig_loopback =-7571;
24479: waveform_sig_loopback =-3274;
24480: waveform_sig_loopback =-6678;
24481: waveform_sig_loopback =-6908;
24482: waveform_sig_loopback =-7321;
24483: waveform_sig_loopback =-5452;
24484: waveform_sig_loopback =-4386;
24485: waveform_sig_loopback =-7463;
24486: waveform_sig_loopback =-6630;
24487: waveform_sig_loopback =-5145;
24488: waveform_sig_loopback =-6668;
24489: waveform_sig_loopback =-5100;
24490: waveform_sig_loopback =-7197;
24491: waveform_sig_loopback =-5600;
24492: waveform_sig_loopback =-4996;
24493: waveform_sig_loopback =-7172;
24494: waveform_sig_loopback =-5353;
24495: waveform_sig_loopback =-5781;
24496: waveform_sig_loopback =-5974;
24497: waveform_sig_loopback =-6271;
24498: waveform_sig_loopback =-4774;
24499: waveform_sig_loopback =-6552;
24500: waveform_sig_loopback =-6013;
24501: waveform_sig_loopback =-4913;
24502: waveform_sig_loopback =-5848;
24503: waveform_sig_loopback =-6201;
24504: waveform_sig_loopback =-5528;
24505: waveform_sig_loopback =-4523;
24506: waveform_sig_loopback =-6781;
24507: waveform_sig_loopback =-5528;
24508: waveform_sig_loopback =-4147;
24509: waveform_sig_loopback =-6511;
24510: waveform_sig_loopback =-6055;
24511: waveform_sig_loopback =-4012;
24512: waveform_sig_loopback =-5483;
24513: waveform_sig_loopback =-6616;
24514: waveform_sig_loopback =-4607;
24515: waveform_sig_loopback =-4486;
24516: waveform_sig_loopback =-6389;
24517: waveform_sig_loopback =-3217;
24518: waveform_sig_loopback =-7503;
24519: waveform_sig_loopback =-6266;
24520: waveform_sig_loopback =-2305;
24521: waveform_sig_loopback =-5405;
24522: waveform_sig_loopback =-5861;
24523: waveform_sig_loopback =-6154;
24524: waveform_sig_loopback =-3993;
24525: waveform_sig_loopback =-3393;
24526: waveform_sig_loopback =-6341;
24527: waveform_sig_loopback =-5155;
24528: waveform_sig_loopback =-4169;
24529: waveform_sig_loopback =-5317;
24530: waveform_sig_loopback =-3832;
24531: waveform_sig_loopback =-6160;
24532: waveform_sig_loopback =-3904;
24533: waveform_sig_loopback =-4073;
24534: waveform_sig_loopback =-5866;
24535: waveform_sig_loopback =-3774;
24536: waveform_sig_loopback =-4858;
24537: waveform_sig_loopback =-4446;
24538: waveform_sig_loopback =-4895;
24539: waveform_sig_loopback =-3682;
24540: waveform_sig_loopback =-4819;
24541: waveform_sig_loopback =-4854;
24542: waveform_sig_loopback =-3631;
24543: waveform_sig_loopback =-4307;
24544: waveform_sig_loopback =-5036;
24545: waveform_sig_loopback =-3652;
24546: waveform_sig_loopback =-3537;
24547: waveform_sig_loopback =-5581;
24548: waveform_sig_loopback =-3645;
24549: waveform_sig_loopback =-2974;
24550: waveform_sig_loopback =-5233;
24551: waveform_sig_loopback =-4503;
24552: waveform_sig_loopback =-2581;
24553: waveform_sig_loopback =-4004;
24554: waveform_sig_loopback =-5215;
24555: waveform_sig_loopback =-3157;
24556: waveform_sig_loopback =-2899;
24557: waveform_sig_loopback =-4931;
24558: waveform_sig_loopback =-1853;
24559: waveform_sig_loopback =-6038;
24560: waveform_sig_loopback =-4497;
24561: waveform_sig_loopback =-914;
24562: waveform_sig_loopback =-3889;
24563: waveform_sig_loopback =-4497;
24564: waveform_sig_loopback =-4472;
24565: waveform_sig_loopback =-2323;
24566: waveform_sig_loopback =-2266;
24567: waveform_sig_loopback =-4537;
24568: waveform_sig_loopback =-3575;
24569: waveform_sig_loopback =-2811;
24570: waveform_sig_loopback =-3396;
24571: waveform_sig_loopback =-2679;
24572: waveform_sig_loopback =-4367;
24573: waveform_sig_loopback =-2147;
24574: waveform_sig_loopback =-2992;
24575: waveform_sig_loopback =-3732;
24576: waveform_sig_loopback =-2451;
24577: waveform_sig_loopback =-3266;
24578: waveform_sig_loopback =-2572;
24579: waveform_sig_loopback =-3678;
24580: waveform_sig_loopback =-1634;
24581: waveform_sig_loopback =-3464;
24582: waveform_sig_loopback =-3299;
24583: waveform_sig_loopback =-1643;
24584: waveform_sig_loopback =-3045;
24585: waveform_sig_loopback =-3254;
24586: waveform_sig_loopback =-1914;
24587: waveform_sig_loopback =-2060;
24588: waveform_sig_loopback =-3815;
24589: waveform_sig_loopback =-1952;
24590: waveform_sig_loopback =-1319;
24591: waveform_sig_loopback =-3665;
24592: waveform_sig_loopback =-2595;
24593: waveform_sig_loopback =-1005;
24594: waveform_sig_loopback =-2330;
24595: waveform_sig_loopback =-3414;
24596: waveform_sig_loopback =-1590;
24597: waveform_sig_loopback =-883;
24598: waveform_sig_loopback =-3406;
24599: waveform_sig_loopback =-111;
24600: waveform_sig_loopback =-4175;
24601: waveform_sig_loopback =-3020;
24602: waveform_sig_loopback =1215;
24603: waveform_sig_loopback =-2371;
24604: waveform_sig_loopback =-2968;
24605: waveform_sig_loopback =-2134;
24606: waveform_sig_loopback =-1081;
24607: waveform_sig_loopback =-243;
24608: waveform_sig_loopback =-2732;
24609: waveform_sig_loopback =-2146;
24610: waveform_sig_loopback =-608;
24611: waveform_sig_loopback =-1887;
24612: waveform_sig_loopback =-873;
24613: waveform_sig_loopback =-2312;
24614: waveform_sig_loopback =-638;
24615: waveform_sig_loopback =-1026;
24616: waveform_sig_loopback =-1895;
24617: waveform_sig_loopback =-826;
24618: waveform_sig_loopback =-1218;
24619: waveform_sig_loopback =-1001;
24620: waveform_sig_loopback =-1719;
24621: waveform_sig_loopback =268;
24622: waveform_sig_loopback =-1799;
24623: waveform_sig_loopback =-1354;
24624: waveform_sig_loopback =248;
24625: waveform_sig_loopback =-1283;
24626: waveform_sig_loopback =-1480;
24627: waveform_sig_loopback =244;
24628: waveform_sig_loopback =-547;
24629: waveform_sig_loopback =-1801;
24630: waveform_sig_loopback =89;
24631: waveform_sig_loopback =154;
24632: waveform_sig_loopback =-1390;
24633: waveform_sig_loopback =-978;
24634: waveform_sig_loopback =918;
24635: waveform_sig_loopback =-208;
24636: waveform_sig_loopback =-2054;
24637: waveform_sig_loopback =839;
24638: waveform_sig_loopback =671;
24639: waveform_sig_loopback =-1712;
24640: waveform_sig_loopback =2296;
24641: waveform_sig_loopback =-2998;
24642: waveform_sig_loopback =-642;
24643: waveform_sig_loopback =3146;
24644: waveform_sig_loopback =-1048;
24645: waveform_sig_loopback =-606;
24646: waveform_sig_loopback =-492;
24647: waveform_sig_loopback =805;
24648: waveform_sig_loopback =1903;
24649: waveform_sig_loopback =-1320;
24650: waveform_sig_loopback =115;
24651: waveform_sig_loopback =1257;
24652: waveform_sig_loopback =-248;
24653: waveform_sig_loopback =1255;
24654: waveform_sig_loopback =-580;
24655: waveform_sig_loopback =1259;
24656: waveform_sig_loopback =950;
24657: waveform_sig_loopback =-123;
24658: waveform_sig_loopback =1108;
24659: waveform_sig_loopback =769;
24660: waveform_sig_loopback =745;
24661: waveform_sig_loopback =221;
24662: waveform_sig_loopback =2304;
24663: waveform_sig_loopback =-211;
24664: waveform_sig_loopback =818;
24665: waveform_sig_loopback =2174;
24666: waveform_sig_loopback =285;
24667: waveform_sig_loopback =856;
24668: waveform_sig_loopback =1882;
24669: waveform_sig_loopback =1264;
24670: waveform_sig_loopback =435;
24671: waveform_sig_loopback =1582;
24672: waveform_sig_loopback =2351;
24673: waveform_sig_loopback =381;
24674: waveform_sig_loopback =707;
24675: waveform_sig_loopback =3308;
24676: waveform_sig_loopback =1121;
24677: waveform_sig_loopback =-48;
24678: waveform_sig_loopback =3174;
24679: waveform_sig_loopback =1891;
24680: waveform_sig_loopback =703;
24681: waveform_sig_loopback =3989;
24682: waveform_sig_loopback =-1510;
24683: waveform_sig_loopback =2022;
24684: waveform_sig_loopback =4414;
24685: waveform_sig_loopback =1033;
24686: waveform_sig_loopback =1438;
24687: waveform_sig_loopback =970;
24688: waveform_sig_loopback =3209;
24689: waveform_sig_loopback =3531;
24690: waveform_sig_loopback =406;
24691: waveform_sig_loopback =2270;
24692: waveform_sig_loopback =2863;
24693: waveform_sig_loopback =1786;
24694: waveform_sig_loopback =3114;
24695: waveform_sig_loopback =1103;
24696: waveform_sig_loopback =3277;
24697: waveform_sig_loopback =2820;
24698: waveform_sig_loopback =1591;
24699: waveform_sig_loopback =2982;
24700: waveform_sig_loopback =2727;
24701: waveform_sig_loopback =2213;
24702: waveform_sig_loopback =2456;
24703: waveform_sig_loopback =3903;
24704: waveform_sig_loopback =1317;
24705: waveform_sig_loopback =3248;
24706: waveform_sig_loopback =3345;
24707: waveform_sig_loopback =2407;
24708: waveform_sig_loopback =2666;
24709: waveform_sig_loopback =3342;
24710: waveform_sig_loopback =3596;
24711: waveform_sig_loopback =1628;
24712: waveform_sig_loopback =3711;
24713: waveform_sig_loopback =4262;
24714: waveform_sig_loopback =1654;
24715: waveform_sig_loopback =3000;
24716: waveform_sig_loopback =4861;
24717: waveform_sig_loopback =2800;
24718: waveform_sig_loopback =1937;
24719: waveform_sig_loopback =4799;
24720: waveform_sig_loopback =3621;
24721: waveform_sig_loopback =2714;
24722: waveform_sig_loopback =5535;
24723: waveform_sig_loopback =142;
24724: waveform_sig_loopback =4180;
24725: waveform_sig_loopback =5859;
24726: waveform_sig_loopback =2882;
24727: waveform_sig_loopback =3099;
24728: waveform_sig_loopback =2608;
24729: waveform_sig_loopback =5282;
24730: waveform_sig_loopback =4875;
24731: waveform_sig_loopback =2090;
24732: waveform_sig_loopback =4284;
24733: waveform_sig_loopback =4161;
24734: waveform_sig_loopback =3747;
24735: waveform_sig_loopback =4696;
24736: waveform_sig_loopback =2597;
24737: waveform_sig_loopback =5331;
24738: waveform_sig_loopback =4128;
24739: waveform_sig_loopback =3299;
24740: waveform_sig_loopback =4898;
24741: waveform_sig_loopback =4060;
24742: waveform_sig_loopback =4030;
24743: waveform_sig_loopback =4247;
24744: waveform_sig_loopback =5247;
24745: waveform_sig_loopback =3286;
24746: waveform_sig_loopback =4694;
24747: waveform_sig_loopback =4868;
24748: waveform_sig_loopback =4316;
24749: waveform_sig_loopback =3937;
24750: waveform_sig_loopback =5219;
24751: waveform_sig_loopback =5143;
24752: waveform_sig_loopback =2960;
24753: waveform_sig_loopback =5731;
24754: waveform_sig_loopback =5596;
24755: waveform_sig_loopback =3076;
24756: waveform_sig_loopback =4954;
24757: waveform_sig_loopback =6105;
24758: waveform_sig_loopback =4405;
24759: waveform_sig_loopback =3679;
24760: waveform_sig_loopback =6147;
24761: waveform_sig_loopback =5256;
24762: waveform_sig_loopback =4255;
24763: waveform_sig_loopback =6821;
24764: waveform_sig_loopback =1795;
24765: waveform_sig_loopback =5711;
24766: waveform_sig_loopback =7273;
24767: waveform_sig_loopback =4436;
24768: waveform_sig_loopback =4313;
24769: waveform_sig_loopback =4377;
24770: waveform_sig_loopback =6733;
24771: waveform_sig_loopback =5999;
24772: waveform_sig_loopback =3865;
24773: waveform_sig_loopback =5670;
24774: waveform_sig_loopback =5416;
24775: waveform_sig_loopback =5469;
24776: waveform_sig_loopback =5796;
24777: waveform_sig_loopback =4208;
24778: waveform_sig_loopback =6837;
24779: waveform_sig_loopback =5129;
24780: waveform_sig_loopback =5083;
24781: waveform_sig_loopback =6111;
24782: waveform_sig_loopback =5313;
24783: waveform_sig_loopback =5650;
24784: waveform_sig_loopback =5358;
24785: waveform_sig_loopback =6619;
24786: waveform_sig_loopback =4751;
24787: waveform_sig_loopback =5743;
24788: waveform_sig_loopback =6485;
24789: waveform_sig_loopback =5471;
24790: waveform_sig_loopback =5055;
24791: waveform_sig_loopback =6859;
24792: waveform_sig_loopback =5955;
24793: waveform_sig_loopback =4463;
24794: waveform_sig_loopback =7168;
24795: waveform_sig_loopback =6379;
24796: waveform_sig_loopback =4588;
24797: waveform_sig_loopback =6237;
24798: waveform_sig_loopback =7140;
24799: waveform_sig_loopback =5741;
24800: waveform_sig_loopback =4776;
24801: waveform_sig_loopback =7412;
24802: waveform_sig_loopback =6468;
24803: waveform_sig_loopback =5320;
24804: waveform_sig_loopback =8067;
24805: waveform_sig_loopback =2894;
24806: waveform_sig_loopback =6871;
24807: waveform_sig_loopback =8561;
24808: waveform_sig_loopback =5404;
24809: waveform_sig_loopback =5254;
24810: waveform_sig_loopback =5901;
24811: waveform_sig_loopback =7618;
24812: waveform_sig_loopback =7172;
24813: waveform_sig_loopback =5005;
24814: waveform_sig_loopback =6576;
24815: waveform_sig_loopback =6716;
24816: waveform_sig_loopback =6469;
24817: waveform_sig_loopback =6665;
24818: waveform_sig_loopback =5531;
24819: waveform_sig_loopback =7706;
24820: waveform_sig_loopback =6116;
24821: waveform_sig_loopback =6369;
24822: waveform_sig_loopback =6762;
24823: waveform_sig_loopback =6565;
24824: waveform_sig_loopback =6626;
24825: waveform_sig_loopback =6123;
24826: waveform_sig_loopback =7956;
24827: waveform_sig_loopback =5401;
24828: waveform_sig_loopback =6828;
24829: waveform_sig_loopback =7631;
24830: waveform_sig_loopback =5996;
24831: waveform_sig_loopback =6358;
24832: waveform_sig_loopback =7823;
24833: waveform_sig_loopback =6522;
24834: waveform_sig_loopback =5812;
24835: waveform_sig_loopback =7839;
24836: waveform_sig_loopback =7229;
24837: waveform_sig_loopback =5652;
24838: waveform_sig_loopback =6833;
24839: waveform_sig_loopback =8176;
24840: waveform_sig_loopback =6426;
24841: waveform_sig_loopback =5483;
24842: waveform_sig_loopback =8539;
24843: waveform_sig_loopback =6943;
24844: waveform_sig_loopback =6243;
24845: waveform_sig_loopback =8876;
24846: waveform_sig_loopback =3366;
24847: waveform_sig_loopback =7916;
24848: waveform_sig_loopback =9249;
24849: waveform_sig_loopback =5842;
24850: waveform_sig_loopback =6187;
24851: waveform_sig_loopback =6428;
24852: waveform_sig_loopback =8216;
24853: waveform_sig_loopback =8072;
24854: waveform_sig_loopback =5437;
24855: waveform_sig_loopback =7046;
24856: waveform_sig_loopback =7623;
24857: waveform_sig_loopback =6991;
24858: waveform_sig_loopback =7306;
24859: waveform_sig_loopback =6148;
24860: waveform_sig_loopback =7976;
24861: waveform_sig_loopback =7194;
24862: waveform_sig_loopback =6592;
24863: waveform_sig_loopback =7188;
24864: waveform_sig_loopback =7506;
24865: waveform_sig_loopback =6610;
24866: waveform_sig_loopback =7074;
24867: waveform_sig_loopback =8218;
24868: waveform_sig_loopback =5679;
24869: waveform_sig_loopback =7776;
24870: waveform_sig_loopback =7706;
24871: waveform_sig_loopback =6499;
24872: waveform_sig_loopback =6961;
24873: waveform_sig_loopback =8060;
24874: waveform_sig_loopback =6982;
24875: waveform_sig_loopback =6134;
24876: waveform_sig_loopback =8184;
24877: waveform_sig_loopback =7691;
24878: waveform_sig_loopback =5922;
24879: waveform_sig_loopback =7163;
24880: waveform_sig_loopback =8714;
24881: waveform_sig_loopback =6579;
24882: waveform_sig_loopback =5750;
24883: waveform_sig_loopback =9133;
24884: waveform_sig_loopback =6816;
24885: waveform_sig_loopback =6828;
24886: waveform_sig_loopback =9079;
24887: waveform_sig_loopback =3290;
24888: waveform_sig_loopback =8846;
24889: waveform_sig_loopback =9112;
24890: waveform_sig_loopback =5960;
24891: waveform_sig_loopback =6727;
24892: waveform_sig_loopback =6456;
24893: waveform_sig_loopback =8631;
24894: waveform_sig_loopback =8118;
24895: waveform_sig_loopback =5287;
24896: waveform_sig_loopback =7941;
24897: waveform_sig_loopback =7347;
24898: waveform_sig_loopback =6961;
24899: waveform_sig_loopback =7773;
24900: waveform_sig_loopback =5937;
24901: waveform_sig_loopback =8460;
24902: waveform_sig_loopback =6987;
24903: waveform_sig_loopback =6520;
24904: waveform_sig_loopback =7731;
24905: waveform_sig_loopback =7238;
24906: waveform_sig_loopback =6634;
24907: waveform_sig_loopback =7338;
24908: waveform_sig_loopback =8011;
24909: waveform_sig_loopback =5845;
24910: waveform_sig_loopback =7729;
24911: waveform_sig_loopback =7514;
24912: waveform_sig_loopback =6663;
24913: waveform_sig_loopback =6846;
24914: waveform_sig_loopback =7899;
24915: waveform_sig_loopback =7037;
24916: waveform_sig_loopback =6085;
24917: waveform_sig_loopback =7995;
24918: waveform_sig_loopback =7681;
24919: waveform_sig_loopback =5643;
24920: waveform_sig_loopback =7223;
24921: waveform_sig_loopback =8645;
24922: waveform_sig_loopback =5951;
24923: waveform_sig_loopback =6113;
24924: waveform_sig_loopback =8855;
24925: waveform_sig_loopback =6261;
24926: waveform_sig_loopback =7295;
24927: waveform_sig_loopback =8266;
24928: waveform_sig_loopback =3254;
24929: waveform_sig_loopback =8920;
24930: waveform_sig_loopback =8335;
24931: waveform_sig_loopback =6216;
24932: waveform_sig_loopback =6128;
24933: waveform_sig_loopback =6179;
24934: waveform_sig_loopback =8796;
24935: waveform_sig_loopback =7262;
24936: waveform_sig_loopback =5196;
24937: waveform_sig_loopback =7725;
24938: waveform_sig_loopback =6619;
24939: waveform_sig_loopback =7100;
24940: waveform_sig_loopback =7052;
24941: waveform_sig_loopback =5565;
24942: waveform_sig_loopback =8431;
24943: waveform_sig_loopback =6168;
24944: waveform_sig_loopback =6408;
24945: waveform_sig_loopback =7215;
24946: waveform_sig_loopback =6701;
24947: waveform_sig_loopback =6367;
24948: waveform_sig_loopback =6826;
24949: waveform_sig_loopback =7475;
24950: waveform_sig_loopback =5423;
24951: waveform_sig_loopback =7309;
24952: waveform_sig_loopback =6824;
24953: waveform_sig_loopback =6328;
24954: waveform_sig_loopback =6195;
24955: waveform_sig_loopback =7340;
24956: waveform_sig_loopback =6659;
24957: waveform_sig_loopback =5185;
24958: waveform_sig_loopback =7805;
24959: waveform_sig_loopback =6929;
24960: waveform_sig_loopback =4781;
24961: waveform_sig_loopback =7166;
24962: waveform_sig_loopback =7481;
24963: waveform_sig_loopback =5467;
24964: waveform_sig_loopback =5722;
24965: waveform_sig_loopback =7752;
24966: waveform_sig_loopback =5989;
24967: waveform_sig_loopback =6431;
24968: waveform_sig_loopback =7380;
24969: waveform_sig_loopback =2938;
24970: waveform_sig_loopback =7932;
24971: waveform_sig_loopback =7841;
24972: waveform_sig_loopback =5401;
24973: waveform_sig_loopback =5135;
24974: waveform_sig_loopback =5833;
24975: waveform_sig_loopback =7766;
24976: waveform_sig_loopback =6491;
24977: waveform_sig_loopback =4552;
24978: waveform_sig_loopback =6823;
24979: waveform_sig_loopback =5844;
24980: waveform_sig_loopback =6357;
24981: waveform_sig_loopback =6077;
24982: waveform_sig_loopback =4869;
24983: waveform_sig_loopback =7575;
24984: waveform_sig_loopback =5036;
24985: waveform_sig_loopback =5823;
24986: waveform_sig_loopback =6289;
24987: waveform_sig_loopback =5611;
24988: waveform_sig_loopback =5731;
24989: waveform_sig_loopback =5793;
24990: waveform_sig_loopback =6508;
24991: waveform_sig_loopback =4719;
24992: waveform_sig_loopback =6013;
24993: waveform_sig_loopback =6277;
24994: waveform_sig_loopback =5172;
24995: waveform_sig_loopback =5105;
24996: waveform_sig_loopback =6812;
24997: waveform_sig_loopback =5077;
24998: waveform_sig_loopback =4523;
24999: waveform_sig_loopback =6887;
25000: waveform_sig_loopback =5484;
25001: waveform_sig_loopback =4119;
25002: waveform_sig_loopback =6034;
25003: waveform_sig_loopback =6359;
25004: waveform_sig_loopback =4518;
25005: waveform_sig_loopback =4484;
25006: waveform_sig_loopback =6849;
25007: waveform_sig_loopback =4790;
25008: waveform_sig_loopback =5309;
25009: waveform_sig_loopback =6238;
25010: waveform_sig_loopback =1760;
25011: waveform_sig_loopback =6904;
25012: waveform_sig_loopback =6690;
25013: waveform_sig_loopback =4069;
25014: waveform_sig_loopback =3952;
25015: waveform_sig_loopback =4898;
25016: waveform_sig_loopback =6401;
25017: waveform_sig_loopback =5275;
25018: waveform_sig_loopback =3432;
25019: waveform_sig_loopback =5495;
25020: waveform_sig_loopback =4772;
25021: waveform_sig_loopback =5121;
25022: waveform_sig_loopback =4564;
25023: waveform_sig_loopback =3990;
25024: waveform_sig_loopback =6097;
25025: waveform_sig_loopback =3710;
25026: waveform_sig_loopback =4805;
25027: waveform_sig_loopback =4628;
25028: waveform_sig_loopback =4659;
25029: waveform_sig_loopback =4256;
25030: waveform_sig_loopback =4370;
25031: waveform_sig_loopback =5504;
25032: waveform_sig_loopback =3013;
25033: waveform_sig_loopback =4872;
25034: waveform_sig_loopback =5008;
25035: waveform_sig_loopback =3446;
25036: waveform_sig_loopback =4152;
25037: waveform_sig_loopback =5281;
25038: waveform_sig_loopback =3529;
25039: waveform_sig_loopback =3463;
25040: waveform_sig_loopback =5274;
25041: waveform_sig_loopback =4069;
25042: waveform_sig_loopback =2788;
25043: waveform_sig_loopback =4542;
25044: waveform_sig_loopback =5001;
25045: waveform_sig_loopback =2996;
25046: waveform_sig_loopback =3018;
25047: waveform_sig_loopback =5582;
25048: waveform_sig_loopback =3117;
25049: waveform_sig_loopback =3937;
25050: waveform_sig_loopback =4741;
25051: waveform_sig_loopback =145;
25052: waveform_sig_loopback =5650;
25053: waveform_sig_loopback =5156;
25054: waveform_sig_loopback =2312;
25055: waveform_sig_loopback =2618;
25056: waveform_sig_loopback =3434;
25057: waveform_sig_loopback =4709;
25058: waveform_sig_loopback =3923;
25059: waveform_sig_loopback =1680;
25060: waveform_sig_loopback =4012;
25061: waveform_sig_loopback =3387;
25062: waveform_sig_loopback =3252;
25063: waveform_sig_loopback =3263;
25064: waveform_sig_loopback =2422;
25065: waveform_sig_loopback =4291;
25066: waveform_sig_loopback =2476;
25067: waveform_sig_loopback =2901;
25068: waveform_sig_loopback =3126;
25069: waveform_sig_loopback =3161;
25070: waveform_sig_loopback =2304;
25071: waveform_sig_loopback =3165;
25072: waveform_sig_loopback =3569;
25073: waveform_sig_loopback =1367;
25074: waveform_sig_loopback =3482;
25075: waveform_sig_loopback =3108;
25076: waveform_sig_loopback =1864;
25077: waveform_sig_loopback =2582;
25078: waveform_sig_loopback =3521;
25079: waveform_sig_loopback =1788;
25080: waveform_sig_loopback =1931;
25081: waveform_sig_loopback =3443;
25082: waveform_sig_loopback =2425;
25083: waveform_sig_loopback =1153;
25084: waveform_sig_loopback =2705;
25085: waveform_sig_loopback =3525;
25086: waveform_sig_loopback =1037;
25087: waveform_sig_loopback =1335;
25088: waveform_sig_loopback =4174;
25089: waveform_sig_loopback =891;
25090: waveform_sig_loopback =2666;
25091: waveform_sig_loopback =2792;
25092: waveform_sig_loopback =-1836;
25093: waveform_sig_loopback =4541;
25094: waveform_sig_loopback =2915;
25095: waveform_sig_loopback =584;
25096: waveform_sig_loopback =1170;
25097: waveform_sig_loopback =1295;
25098: waveform_sig_loopback =3310;
25099: waveform_sig_loopback =1938;
25100: waveform_sig_loopback =-253;
25101: waveform_sig_loopback =2644;
25102: waveform_sig_loopback =1189;
25103: waveform_sig_loopback =1625;
25104: waveform_sig_loopback =1460;
25105: waveform_sig_loopback =463;
25106: waveform_sig_loopback =2678;
25107: waveform_sig_loopback =538;
25108: waveform_sig_loopback =1090;
25109: waveform_sig_loopback =1412;
25110: waveform_sig_loopback =1271;
25111: waveform_sig_loopback =396;
25112: waveform_sig_loopback =1531;
25113: waveform_sig_loopback =1586;
25114: waveform_sig_loopback =-520;
25115: waveform_sig_loopback =1904;
25116: waveform_sig_loopback =1018;
25117: waveform_sig_loopback =23;
25118: waveform_sig_loopback =978;
25119: waveform_sig_loopback =1308;
25120: waveform_sig_loopback =260;
25121: waveform_sig_loopback =-96;
25122: waveform_sig_loopback =1586;
25123: waveform_sig_loopback =779;
25124: waveform_sig_loopback =-1119;
25125: waveform_sig_loopback =1271;
25126: waveform_sig_loopback =1530;
25127: waveform_sig_loopback =-1092;
25128: waveform_sig_loopback =-43;
25129: waveform_sig_loopback =2008;
25130: waveform_sig_loopback =-1037;
25131: waveform_sig_loopback =1110;
25132: waveform_sig_loopback =441;
25133: waveform_sig_loopback =-3395;
25134: waveform_sig_loopback =2740;
25135: waveform_sig_loopback =668;
25136: waveform_sig_loopback =-935;
25137: waveform_sig_loopback =-964;
25138: waveform_sig_loopback =-539;
25139: waveform_sig_loopback =1709;
25140: waveform_sig_loopback =-379;
25141: waveform_sig_loopback =-1934;
25142: waveform_sig_loopback =808;
25143: waveform_sig_loopback =-862;
25144: waveform_sig_loopback =60;
25145: waveform_sig_loopback =-725;
25146: waveform_sig_loopback =-1387;
25147: waveform_sig_loopback =1002;
25148: waveform_sig_loopback =-1532;
25149: waveform_sig_loopback =-724;
25150: waveform_sig_loopback =-437;
25151: waveform_sig_loopback =-707;
25152: waveform_sig_loopback =-1376;
25153: waveform_sig_loopback =-191;
25154: waveform_sig_loopback =-678;
25155: waveform_sig_loopback =-2117;
25156: waveform_sig_loopback =72;
25157: waveform_sig_loopback =-1177;
25158: waveform_sig_loopback =-1430;
25159: waveform_sig_loopback =-1287;
25160: waveform_sig_loopback =-308;
25161: waveform_sig_loopback =-1603;
25162: waveform_sig_loopback =-2315;
25163: waveform_sig_loopback =260;
25164: waveform_sig_loopback =-1517;
25165: waveform_sig_loopback =-2975;
25166: waveform_sig_loopback =-281;
25167: waveform_sig_loopback =-737;
25168: waveform_sig_loopback =-2782;
25169: waveform_sig_loopback =-1940;
25170: waveform_sig_loopback =8;
25171: waveform_sig_loopback =-2747;
25172: waveform_sig_loopback =-710;
25173: waveform_sig_loopback =-1760;
25174: waveform_sig_loopback =-4948;
25175: waveform_sig_loopback =912;
25176: waveform_sig_loopback =-1383;
25177: waveform_sig_loopback =-2657;
25178: waveform_sig_loopback =-3022;
25179: waveform_sig_loopback =-2174;
25180: waveform_sig_loopback =-91;
25181: waveform_sig_loopback =-2550;
25182: waveform_sig_loopback =-3466;
25183: waveform_sig_loopback =-1147;
25184: waveform_sig_loopback =-2873;
25185: waveform_sig_loopback =-1513;
25186: waveform_sig_loopback =-2892;
25187: waveform_sig_loopback =-2938;
25188: waveform_sig_loopback =-875;
25189: waveform_sig_loopback =-3718;
25190: waveform_sig_loopback =-2174;
25191: waveform_sig_loopback =-2351;
25192: waveform_sig_loopback =-2757;
25193: waveform_sig_loopback =-2971;
25194: waveform_sig_loopback =-2154;
25195: waveform_sig_loopback =-2616;
25196: waveform_sig_loopback =-3724;
25197: waveform_sig_loopback =-2105;
25198: waveform_sig_loopback =-2731;
25199: waveform_sig_loopback =-3395;
25200: waveform_sig_loopback =-3416;
25201: waveform_sig_loopback =-1716;
25202: waveform_sig_loopback =-3819;
25203: waveform_sig_loopback =-3891;
25204: waveform_sig_loopback =-1638;
25205: waveform_sig_loopback =-3703;
25206: waveform_sig_loopback =-4253;
25207: waveform_sig_loopback =-2208;
25208: waveform_sig_loopback =-2800;
25209: waveform_sig_loopback =-4458;
25210: waveform_sig_loopback =-3565;
25211: waveform_sig_loopback =-1855;
25212: waveform_sig_loopback =-4609;
25213: waveform_sig_loopback =-2434;
25214: waveform_sig_loopback =-3659;
25215: waveform_sig_loopback =-6514;
25216: waveform_sig_loopback =-1056;
25217: waveform_sig_loopback =-2993;
25218: waveform_sig_loopback =-4466;
25219: waveform_sig_loopback =-4949;
25220: waveform_sig_loopback =-3542;
25221: waveform_sig_loopback =-2116;
25222: waveform_sig_loopback =-4262;
25223: waveform_sig_loopback =-4980;
25224: waveform_sig_loopback =-3216;
25225: waveform_sig_loopback =-4266;
25226: waveform_sig_loopback =-3343;
25227: waveform_sig_loopback =-4808;
25228: waveform_sig_loopback =-4241;
25229: waveform_sig_loopback =-2936;
25230: waveform_sig_loopback =-5297;
25231: waveform_sig_loopback =-3776;
25232: waveform_sig_loopback =-4338;
25233: waveform_sig_loopback =-4154;
25234: waveform_sig_loopback =-4756;
25235: waveform_sig_loopback =-3894;
25236: waveform_sig_loopback =-4102;
25237: waveform_sig_loopback =-5458;
25238: waveform_sig_loopback =-3777;
25239: waveform_sig_loopback =-4164;
25240: waveform_sig_loopback =-5317;
25241: waveform_sig_loopback =-4595;
25242: waveform_sig_loopback =-3322;
25243: waveform_sig_loopback =-5885;
25244: waveform_sig_loopback =-4935;
25245: waveform_sig_loopback =-3264;
25246: waveform_sig_loopback =-5440;
25247: waveform_sig_loopback =-5674;
25248: waveform_sig_loopback =-3985;
25249: waveform_sig_loopback =-4044;
25250: waveform_sig_loopback =-6034;
25251: waveform_sig_loopback =-5402;
25252: waveform_sig_loopback =-3017;
25253: waveform_sig_loopback =-6314;
25254: waveform_sig_loopback =-3899;
25255: waveform_sig_loopback =-5209;
25256: waveform_sig_loopback =-8094;
25257: waveform_sig_loopback =-2263;
25258: waveform_sig_loopback =-4594;
25259: waveform_sig_loopback =-6227;
25260: waveform_sig_loopback =-6152;
25261: waveform_sig_loopback =-4932;
25262: waveform_sig_loopback =-3813;
25263: waveform_sig_loopback =-5626;
25264: waveform_sig_loopback =-6477;
25265: waveform_sig_loopback =-4620;
25266: waveform_sig_loopback =-5500;
25267: waveform_sig_loopback =-5059;
25268: waveform_sig_loopback =-6061;
25269: waveform_sig_loopback =-5488;
25270: waveform_sig_loopback =-4642;
25271: waveform_sig_loopback =-6311;
25272: waveform_sig_loopback =-5295;
25273: waveform_sig_loopback =-5751;
25274: waveform_sig_loopback =-5214;
25275: waveform_sig_loopback =-6525;
25276: waveform_sig_loopback =-4940;
25277: waveform_sig_loopback =-5446;
25278: waveform_sig_loopback =-7089;
25279: waveform_sig_loopback =-4699;
25280: waveform_sig_loopback =-5705;
25281: waveform_sig_loopback =-6693;
25282: waveform_sig_loopback =-5570;
25283: waveform_sig_loopback =-5015;
25284: waveform_sig_loopback =-7031;
25285: waveform_sig_loopback =-6041;
25286: waveform_sig_loopback =-4817;
25287: waveform_sig_loopback =-6471;
25288: waveform_sig_loopback =-7032;
25289: waveform_sig_loopback =-5226;
25290: waveform_sig_loopback =-5121;
25291: waveform_sig_loopback =-7579;
25292: waveform_sig_loopback =-6364;
25293: waveform_sig_loopback =-4169;
25294: waveform_sig_loopback =-7800;
25295: waveform_sig_loopback =-4724;
25296: waveform_sig_loopback =-6724;
25297: waveform_sig_loopback =-9188;
25298: waveform_sig_loopback =-3150;
25299: waveform_sig_loopback =-6056;
25300: waveform_sig_loopback =-7358;
25301: waveform_sig_loopback =-7056;
25302: waveform_sig_loopback =-6222;
25303: waveform_sig_loopback =-4769;
25304: waveform_sig_loopback =-6714;
25305: waveform_sig_loopback =-7820;
25306: waveform_sig_loopback =-5375;
25307: waveform_sig_loopback =-6744;
25308: waveform_sig_loopback =-6182;
25309: waveform_sig_loopback =-6856;
25310: waveform_sig_loopback =-6730;
25311: waveform_sig_loopback =-5586;
25312: waveform_sig_loopback =-7218;
25313: waveform_sig_loopback =-6576;
25314: waveform_sig_loopback =-6441;
25315: waveform_sig_loopback =-6315;
25316: waveform_sig_loopback =-7651;
25317: waveform_sig_loopback =-5415;
25318: waveform_sig_loopback =-6932;
25319: waveform_sig_loopback =-7741;
25320: waveform_sig_loopback =-5433;
25321: waveform_sig_loopback =-7074;
25322: waveform_sig_loopback =-7163;
25323: waveform_sig_loopback =-6624;
25324: waveform_sig_loopback =-5951;
25325: waveform_sig_loopback =-7672;
25326: waveform_sig_loopback =-7098;
25327: waveform_sig_loopback =-5523;
25328: waveform_sig_loopback =-7359;
25329: waveform_sig_loopback =-7925;
25330: waveform_sig_loopback =-5874;
25331: waveform_sig_loopback =-6035;
25332: waveform_sig_loopback =-8504;
25333: waveform_sig_loopback =-6956;
25334: waveform_sig_loopback =-5033;
25335: waveform_sig_loopback =-8762;
25336: waveform_sig_loopback =-5075;
25337: waveform_sig_loopback =-7906;
25338: waveform_sig_loopback =-9742;
25339: waveform_sig_loopback =-3519;
25340: waveform_sig_loopback =-7274;
25341: waveform_sig_loopback =-7801;
25342: waveform_sig_loopback =-7718;
25343: waveform_sig_loopback =-7163;
25344: waveform_sig_loopback =-4963;
25345: waveform_sig_loopback =-7852;
25346: waveform_sig_loopback =-8296;
25347: waveform_sig_loopback =-5694;
25348: waveform_sig_loopback =-7923;
25349: waveform_sig_loopback =-6323;
25350: waveform_sig_loopback =-7687;
25351: waveform_sig_loopback =-7450;
25352: waveform_sig_loopback =-5769;
25353: waveform_sig_loopback =-8290;
25354: waveform_sig_loopback =-6883;
25355: waveform_sig_loopback =-6861;
25356: waveform_sig_loopback =-7241;
25357: waveform_sig_loopback =-7748;
25358: waveform_sig_loopback =-6126;
25359: waveform_sig_loopback =-7498;
25360: waveform_sig_loopback =-7933;
25361: waveform_sig_loopback =-6170;
25362: waveform_sig_loopback =-7397;
25363: waveform_sig_loopback =-7637;
25364: waveform_sig_loopback =-6996;
25365: waveform_sig_loopback =-6426;
25366: waveform_sig_loopback =-8115;
25367: waveform_sig_loopback =-7501;
25368: waveform_sig_loopback =-5871;
25369: waveform_sig_loopback =-7751;
25370: waveform_sig_loopback =-8467;
25371: waveform_sig_loopback =-5880;
25372: waveform_sig_loopback =-6596;
25373: waveform_sig_loopback =-8982;
25374: waveform_sig_loopback =-6757;
25375: waveform_sig_loopback =-5849;
25376: waveform_sig_loopback =-8768;
25377: waveform_sig_loopback =-5184;
25378: waveform_sig_loopback =-8877;
25379: waveform_sig_loopback =-9196;
25380: waveform_sig_loopback =-4169;
25381: waveform_sig_loopback =-7574;
25382: waveform_sig_loopback =-7647;
25383: waveform_sig_loopback =-8555;
25384: waveform_sig_loopback =-6720;
25385: waveform_sig_loopback =-5351;
25386: waveform_sig_loopback =-8395;
25387: waveform_sig_loopback =-7847;
25388: waveform_sig_loopback =-6370;
25389: waveform_sig_loopback =-7809;
25390: waveform_sig_loopback =-6311;
25391: waveform_sig_loopback =-8318;
25392: waveform_sig_loopback =-7015;
25393: waveform_sig_loopback =-6132;
25394: waveform_sig_loopback =-8482;
25395: waveform_sig_loopback =-6655;
25396: waveform_sig_loopback =-7179;
25397: waveform_sig_loopback =-7119;
25398: waveform_sig_loopback =-7837;
25399: waveform_sig_loopback =-6281;
25400: waveform_sig_loopback =-7446;
25401: waveform_sig_loopback =-7816;
25402: waveform_sig_loopback =-6227;
25403: waveform_sig_loopback =-7366;
25404: waveform_sig_loopback =-7679;
25405: waveform_sig_loopback =-7137;
25406: waveform_sig_loopback =-5990;
25407: waveform_sig_loopback =-8123;
25408: waveform_sig_loopback =-7606;
25409: waveform_sig_loopback =-5607;
25410: waveform_sig_loopback =-7945;
25411: waveform_sig_loopback =-7909;
25412: waveform_sig_loopback =-5765;
25413: waveform_sig_loopback =-6999;
25414: waveform_sig_loopback =-8205;
25415: waveform_sig_loopback =-6770;
25416: waveform_sig_loopback =-5834;
25417: waveform_sig_loopback =-8192;
25418: waveform_sig_loopback =-5404;
25419: waveform_sig_loopback =-8477;
25420: waveform_sig_loopback =-8919;
25421: waveform_sig_loopback =-4143;
25422: waveform_sig_loopback =-6795;
25423: waveform_sig_loopback =-8001;
25424: waveform_sig_loopback =-8113;
25425: waveform_sig_loopback =-6085;
25426: waveform_sig_loopback =-5477;
25427: waveform_sig_loopback =-7757;
25428: waveform_sig_loopback =-7782;
25429: waveform_sig_loopback =-6034;
25430: waveform_sig_loopback =-7126;
25431: waveform_sig_loopback =-6274;
25432: waveform_sig_loopback =-7848;
25433: waveform_sig_loopback =-6509;
25434: waveform_sig_loopback =-5955;
25435: waveform_sig_loopback =-7918;
25436: waveform_sig_loopback =-6292;
25437: waveform_sig_loopback =-6782;
25438: waveform_sig_loopback =-6714;
25439: waveform_sig_loopback =-7366;
25440: waveform_sig_loopback =-5839;
25441: waveform_sig_loopback =-6915;
25442: waveform_sig_loopback =-7324;
25443: waveform_sig_loopback =-5985;
25444: waveform_sig_loopback =-6458;
25445: waveform_sig_loopback =-7446;
25446: waveform_sig_loopback =-6344;
25447: waveform_sig_loopback =-5566;
25448: waveform_sig_loopback =-8101;
25449: waveform_sig_loopback =-6207;
25450: waveform_sig_loopback =-5449;
25451: waveform_sig_loopback =-7505;
25452: waveform_sig_loopback =-7024;
25453: waveform_sig_loopback =-5510;
25454: waveform_sig_loopback =-5960;
25455: waveform_sig_loopback =-7926;
25456: waveform_sig_loopback =-6189;
25457: waveform_sig_loopback =-4811;
25458: waveform_sig_loopback =-8014;
25459: waveform_sig_loopback =-4422;
25460: waveform_sig_loopback =-7934;
25461: waveform_sig_loopback =-8255;
25462: waveform_sig_loopback =-3139;
25463: waveform_sig_loopback =-6485;
25464: waveform_sig_loopback =-7226;
25465: waveform_sig_loopback =-6977;
25466: waveform_sig_loopback =-5650;
25467: waveform_sig_loopback =-4651;
25468: waveform_sig_loopback =-6976;
25469: waveform_sig_loopback =-6968;
25470: waveform_sig_loopback =-5121;
25471: waveform_sig_loopback =-6482;
25472: waveform_sig_loopback =-5424;
25473: waveform_sig_loopback =-6892;
25474: waveform_sig_loopback =-5639;
25475: waveform_sig_loopback =-5228;
25476: waveform_sig_loopback =-6883;
25477: waveform_sig_loopback =-5425;
25478: waveform_sig_loopback =-5989;
25479: waveform_sig_loopback =-5610;
25480: waveform_sig_loopback =-6610;
25481: waveform_sig_loopback =-4751;
25482: waveform_sig_loopback =-5985;
25483: waveform_sig_loopback =-6714;
25484: waveform_sig_loopback =-4517;
25485: waveform_sig_loopback =-5892;
25486: waveform_sig_loopback =-6477;
25487: waveform_sig_loopback =-4868;
25488: waveform_sig_loopback =-5193;
25489: waveform_sig_loopback =-6603;
25490: waveform_sig_loopback =-5348;
25491: waveform_sig_loopback =-4514;
25492: waveform_sig_loopback =-6116;
25493: waveform_sig_loopback =-6320;
25494: waveform_sig_loopback =-4185;
25495: waveform_sig_loopback =-4997;
25496: waveform_sig_loopback =-6944;
25497: waveform_sig_loopback =-4692;
25498: waveform_sig_loopback =-4006;
25499: waveform_sig_loopback =-6837;
25500: waveform_sig_loopback =-3092;
25501: waveform_sig_loopback =-7100;
25502: waveform_sig_loopback =-6823;
25503: waveform_sig_loopback =-1879;
25504: waveform_sig_loopback =-5570;
25505: waveform_sig_loopback =-5968;
25506: waveform_sig_loopback =-5683;
25507: waveform_sig_loopback =-4519;
25508: waveform_sig_loopback =-3265;
25509: waveform_sig_loopback =-5952;
25510: waveform_sig_loopback =-5694;
25511: waveform_sig_loopback =-3792;
25512: waveform_sig_loopback =-5402;
25513: waveform_sig_loopback =-4089;
25514: waveform_sig_loopback =-5620;
25515: waveform_sig_loopback =-4409;
25516: waveform_sig_loopback =-3914;
25517: waveform_sig_loopback =-5525;
25518: waveform_sig_loopback =-4271;
25519: waveform_sig_loopback =-4479;
25520: waveform_sig_loopback =-4424;
25521: waveform_sig_loopback =-5332;
25522: waveform_sig_loopback =-3078;
25523: waveform_sig_loopback =-5075;
25524: waveform_sig_loopback =-5022;
25525: waveform_sig_loopback =-3114;
25526: waveform_sig_loopback =-4803;
25527: waveform_sig_loopback =-4683;
25528: waveform_sig_loopback =-3766;
25529: waveform_sig_loopback =-3742;
25530: waveform_sig_loopback =-5020;
25531: waveform_sig_loopback =-4168;
25532: waveform_sig_loopback =-2848;
25533: waveform_sig_loopback =-4863;
25534: waveform_sig_loopback =-4903;
25535: waveform_sig_loopback =-2450;
25536: waveform_sig_loopback =-3826;
25537: waveform_sig_loopback =-5435;
25538: waveform_sig_loopback =-3072;
25539: waveform_sig_loopback =-2727;
25540: waveform_sig_loopback =-5237;
25541: waveform_sig_loopback =-1526;
25542: waveform_sig_loopback =-5987;
25543: waveform_sig_loopback =-4984;
25544: waveform_sig_loopback =-391;
25545: waveform_sig_loopback =-4281;
25546: waveform_sig_loopback =-4249;
25547: waveform_sig_loopback =-4374;
25548: waveform_sig_loopback =-3123;
25549: waveform_sig_loopback =-1398;
25550: waveform_sig_loopback =-4781;
25551: waveform_sig_loopback =-3943;
25552: waveform_sig_loopback =-2419;
25553: waveform_sig_loopback =-3906;
25554: waveform_sig_loopback =-2084;
25555: waveform_sig_loopback =-4455;
25556: waveform_sig_loopback =-2794;
25557: waveform_sig_loopback =-2171;
25558: waveform_sig_loopback =-4077;
25559: waveform_sig_loopback =-2597;
25560: waveform_sig_loopback =-2934;
25561: waveform_sig_loopback =-2984;
25562: waveform_sig_loopback =-3383;
25563: waveform_sig_loopback =-1704;
25564: waveform_sig_loopback =-3631;
25565: waveform_sig_loopback =-3012;
25566: waveform_sig_loopback =-1744;
25567: waveform_sig_loopback =-3132;
25568: waveform_sig_loopback =-3040;
25569: waveform_sig_loopback =-2131;
25570: waveform_sig_loopback =-1959;
25571: waveform_sig_loopback =-3569;
25572: waveform_sig_loopback =-2462;
25573: waveform_sig_loopback =-1004;
25574: waveform_sig_loopback =-3387;
25575: waveform_sig_loopback =-3220;
25576: waveform_sig_loopback =-559;
25577: waveform_sig_loopback =-2398;
25578: waveform_sig_loopback =-3567;
25579: waveform_sig_loopback =-1272;
25580: waveform_sig_loopback =-1362;
25581: waveform_sig_loopback =-3094;
25582: waveform_sig_loopback =20;
25583: waveform_sig_loopback =-4516;
25584: waveform_sig_loopback =-2708;
25585: waveform_sig_loopback =1024;
25586: waveform_sig_loopback =-2409;
25587: waveform_sig_loopback =-2497;
25588: waveform_sig_loopback =-2791;
25589: waveform_sig_loopback =-775;
25590: waveform_sig_loopback =-25;
25591: waveform_sig_loopback =-3180;
25592: waveform_sig_loopback =-1745;
25593: waveform_sig_loopback =-784;
25594: waveform_sig_loopback =-2053;
25595: waveform_sig_loopback =-422;
25596: waveform_sig_loopback =-2826;
25597: waveform_sig_loopback =-523;
25598: waveform_sig_loopback =-651;
25599: waveform_sig_loopback =-2446;
25600: waveform_sig_loopback =-469;
25601: waveform_sig_loopback =-1240;
25602: waveform_sig_loopback =-1181;
25603: waveform_sig_loopback =-1421;
25604: waveform_sig_loopback =-20;
25605: waveform_sig_loopback =-1677;
25606: waveform_sig_loopback =-1127;
25607: waveform_sig_loopback =-204;
25608: waveform_sig_loopback =-945;
25609: waveform_sig_loopback =-1392;
25610: waveform_sig_loopback =-311;
25611: waveform_sig_loopback =63;
25612: waveform_sig_loopback =-1997;
25613: waveform_sig_loopback =-222;
25614: waveform_sig_loopback =669;
25615: waveform_sig_loopback =-1758;
25616: waveform_sig_loopback =-925;
25617: waveform_sig_loopback =1061;
25618: waveform_sig_loopback =-593;
25619: waveform_sig_loopback =-1555;
25620: waveform_sig_loopback =571;
25621: waveform_sig_loopback =500;
25622: waveform_sig_loopback =-1188;
25623: waveform_sig_loopback =1820;
25624: waveform_sig_loopback =-2662;
25625: waveform_sig_loopback =-609;
25626: waveform_sig_loopback =2657;
25627: waveform_sig_loopback =-405;
25628: waveform_sig_loopback =-774;
25629: waveform_sig_loopback =-804;
25630: waveform_sig_loopback =1232;
25631: waveform_sig_loopback =1648;
25632: waveform_sig_loopback =-1198;
25633: waveform_sig_loopback =301;
25634: waveform_sig_loopback =833;
25635: waveform_sig_loopback =173;
25636: waveform_sig_loopback =1316;
25637: waveform_sig_loopback =-996;
25638: waveform_sig_loopback =1739;
25639: waveform_sig_loopback =766;
25640: waveform_sig_loopback =-202;
25641: waveform_sig_loopback =1372;
25642: waveform_sig_loopback =420;
25643: waveform_sig_loopback =1030;
25644: waveform_sig_loopback =223;
25645: waveform_sig_loopback =1965;
25646: waveform_sig_loopback =229;
25647: waveform_sig_loopback =630;
25648: waveform_sig_loopback =1881;
25649: waveform_sig_loopback =824;
25650: waveform_sig_loopback =387;
25651: waveform_sig_loopback =1861;
25652: waveform_sig_loopback =1745;
25653: waveform_sig_loopback =-173;
25654: waveform_sig_loopback =1946;
25655: waveform_sig_loopback =2322;
25656: waveform_sig_loopback =135;
25657: waveform_sig_loopback =1139;
25658: waveform_sig_loopback =2788;
25659: waveform_sig_loopback =1381;
25660: waveform_sig_loopback =305;
25661: waveform_sig_loopback =2465;
25662: waveform_sig_loopback =2425;
25663: waveform_sig_loopback =639;
25664: waveform_sig_loopback =3689;
25665: waveform_sig_loopback =-882;
25666: waveform_sig_loopback =1358;
25667: waveform_sig_loopback =4618;
25668: waveform_sig_loopback =1414;
25669: waveform_sig_loopback =860;
25670: waveform_sig_loopback =1306;
25671: waveform_sig_loopback =3139;
25672: waveform_sig_loopback =3203;
25673: waveform_sig_loopback =895;
25674: waveform_sig_loopback =1945;
25675: waveform_sig_loopback =2792;
25676: waveform_sig_loopback =2108;
25677: waveform_sig_loopback =2748;
25678: waveform_sig_loopback =1255;
25679: waveform_sig_loopback =3377;
25680: waveform_sig_loopback =2466;
25681: waveform_sig_loopback =1932;
25682: waveform_sig_loopback =2924;
25683: waveform_sig_loopback =2497;
25684: waveform_sig_loopback =2751;
25685: waveform_sig_loopback =1963;
25686: waveform_sig_loopback =4023;
25687: waveform_sig_loopback =1818;
25688: waveform_sig_loopback =2535;
25689: waveform_sig_loopback =3771;
25690: waveform_sig_loopback =2470;
25691: waveform_sig_loopback =2334;
25692: waveform_sig_loopback =3719;
25693: waveform_sig_loopback =3356;
25694: waveform_sig_loopback =1707;
25695: waveform_sig_loopback =3872;
25696: waveform_sig_loopback =3915;
25697: waveform_sig_loopback =1938;
25698: waveform_sig_loopback =3080;
25699: waveform_sig_loopback =4382;
25700: waveform_sig_loopback =3254;
25701: waveform_sig_loopback =1854;
25702: waveform_sig_loopback =4363;
25703: waveform_sig_loopback =4257;
25704: waveform_sig_loopback =2028;
25705: waveform_sig_loopback =5773;
25706: waveform_sig_loopback =563;
25707: waveform_sig_loopback =3251;
25708: waveform_sig_loopback =6571;
25709: waveform_sig_loopback =2622;
25710: waveform_sig_loopback =2849;
25711: waveform_sig_loopback =3163;
25712: waveform_sig_loopback =4607;
25713: waveform_sig_loopback =5158;
25714: waveform_sig_loopback =2351;
25715: waveform_sig_loopback =3775;
25716: waveform_sig_loopback =4655;
25717: waveform_sig_loopback =3570;
25718: waveform_sig_loopback =4597;
25719: waveform_sig_loopback =2978;
25720: waveform_sig_loopback =4957;
25721: waveform_sig_loopback =4259;
25722: waveform_sig_loopback =3516;
25723: waveform_sig_loopback =4534;
25724: waveform_sig_loopback =4266;
25725: waveform_sig_loopback =4253;
25726: waveform_sig_loopback =3650;
25727: waveform_sig_loopback =5725;
25728: waveform_sig_loopback =3290;
25729: waveform_sig_loopback =4251;
25730: waveform_sig_loopback =5442;
25731: waveform_sig_loopback =3845;
25732: waveform_sig_loopback =4119;
25733: waveform_sig_loopback =5336;
25734: waveform_sig_loopback =4668;
25735: waveform_sig_loopback =3593;
25736: waveform_sig_loopback =5300;
25737: waveform_sig_loopback =5443;
25738: waveform_sig_loopback =3638;
25739: waveform_sig_loopback =4387;
25740: waveform_sig_loopback =6289;
25741: waveform_sig_loopback =4604;
25742: waveform_sig_loopback =3265;
25743: waveform_sig_loopback =6396;
25744: waveform_sig_loopback =5285;
25745: waveform_sig_loopback =3892;
25746: waveform_sig_loopback =7328;
25747: waveform_sig_loopback =1584;
25748: waveform_sig_loopback =5419;
25749: waveform_sig_loopback =7733;
25750: waveform_sig_loopback =4015;
25751: waveform_sig_loopback =4558;
25752: waveform_sig_loopback =4441;
25753: waveform_sig_loopback =6298;
25754: waveform_sig_loopback =6560;
25755: waveform_sig_loopback =3601;
25756: waveform_sig_loopback =5455;
25757: waveform_sig_loopback =5942;
25758: waveform_sig_loopback =4963;
25759: waveform_sig_loopback =6049;
25760: waveform_sig_loopback =4329;
25761: waveform_sig_loopback =6358;
25762: waveform_sig_loopback =5703;
25763: waveform_sig_loopback =4828;
25764: waveform_sig_loopback =5869;
25765: waveform_sig_loopback =5853;
25766: waveform_sig_loopback =5274;
25767: waveform_sig_loopback =5264;
25768: waveform_sig_loopback =7027;
25769: waveform_sig_loopback =4289;
25770: waveform_sig_loopback =6087;
25771: waveform_sig_loopback =6392;
25772: waveform_sig_loopback =5194;
25773: waveform_sig_loopback =5648;
25774: waveform_sig_loopback =6346;
25775: waveform_sig_loopback =6150;
25776: waveform_sig_loopback =4785;
25777: waveform_sig_loopback =6544;
25778: waveform_sig_loopback =6850;
25779: waveform_sig_loopback =4633;
25780: waveform_sig_loopback =5795;
25781: waveform_sig_loopback =7542;
25782: waveform_sig_loopback =5505;
25783: waveform_sig_loopback =4668;
25784: waveform_sig_loopback =7675;
25785: waveform_sig_loopback =6114;
25786: waveform_sig_loopback =5385;
25787: waveform_sig_loopback =8275;
25788: waveform_sig_loopback =2608;
25789: waveform_sig_loopback =6976;
25790: waveform_sig_loopback =8525;
25791: waveform_sig_loopback =5248;
25792: waveform_sig_loopback =5711;
25793: waveform_sig_loopback =5350;
25794: waveform_sig_loopback =7673;
25795: waveform_sig_loopback =7559;
25796: waveform_sig_loopback =4521;
25797: waveform_sig_loopback =6789;
25798: waveform_sig_loopback =6779;
25799: waveform_sig_loopback =6092;
25800: waveform_sig_loopback =7222;
25801: waveform_sig_loopback =5052;
25802: waveform_sig_loopback =7649;
25803: waveform_sig_loopback =6686;
25804: waveform_sig_loopback =5617;
25805: waveform_sig_loopback =7187;
25806: waveform_sig_loopback =6601;
25807: waveform_sig_loopback =6209;
25808: waveform_sig_loopback =6620;
25809: waveform_sig_loopback =7530;
25810: waveform_sig_loopback =5535;
25811: waveform_sig_loopback =7035;
25812: waveform_sig_loopback =7025;
25813: waveform_sig_loopback =6493;
25814: waveform_sig_loopback =6216;
25815: waveform_sig_loopback =7421;
25816: waveform_sig_loopback =7081;
25817: waveform_sig_loopback =5407;
25818: waveform_sig_loopback =7738;
25819: waveform_sig_loopback =7504;
25820: waveform_sig_loopback =5442;
25821: waveform_sig_loopback =6801;
25822: waveform_sig_loopback =8288;
25823: waveform_sig_loopback =6259;
25824: waveform_sig_loopback =5606;
25825: waveform_sig_loopback =8526;
25826: waveform_sig_loopback =6639;
25827: waveform_sig_loopback =6560;
25828: waveform_sig_loopback =8755;
25829: waveform_sig_loopback =3275;
25830: waveform_sig_loopback =8172;
25831: waveform_sig_loopback =8757;
25832: waveform_sig_loopback =6301;
25833: waveform_sig_loopback =6266;
25834: waveform_sig_loopback =5985;
25835: waveform_sig_loopback =8811;
25836: waveform_sig_loopback =7639;
25837: waveform_sig_loopback =5456;
25838: waveform_sig_loopback =7620;
25839: waveform_sig_loopback =7025;
25840: waveform_sig_loopback =7207;
25841: waveform_sig_loopback =7478;
25842: waveform_sig_loopback =5800;
25843: waveform_sig_loopback =8529;
25844: waveform_sig_loopback =6738;
25845: waveform_sig_loopback =6573;
25846: waveform_sig_loopback =7745;
25847: waveform_sig_loopback =6966;
25848: waveform_sig_loopback =6986;
25849: waveform_sig_loopback =6935;
25850: waveform_sig_loopback =8147;
25851: waveform_sig_loopback =6076;
25852: waveform_sig_loopback =7446;
25853: waveform_sig_loopback =7626;
25854: waveform_sig_loopback =6893;
25855: waveform_sig_loopback =6707;
25856: waveform_sig_loopback =7912;
25857: waveform_sig_loopback =7490;
25858: waveform_sig_loopback =5722;
25859: waveform_sig_loopback =8355;
25860: waveform_sig_loopback =7819;
25861: waveform_sig_loopback =5583;
25862: waveform_sig_loopback =7707;
25863: waveform_sig_loopback =8306;
25864: waveform_sig_loopback =6592;
25865: waveform_sig_loopback =6215;
25866: waveform_sig_loopback =8541;
25867: waveform_sig_loopback =7263;
25868: waveform_sig_loopback =6741;
25869: waveform_sig_loopback =8859;
25870: waveform_sig_loopback =3883;
25871: waveform_sig_loopback =8237;
25872: waveform_sig_loopback =9214;
25873: waveform_sig_loopback =6556;
25874: waveform_sig_loopback =6123;
25875: waveform_sig_loopback =6696;
25876: waveform_sig_loopback =8838;
25877: waveform_sig_loopback =7746;
25878: waveform_sig_loopback =5879;
25879: waveform_sig_loopback =7521;
25880: waveform_sig_loopback =7344;
25881: waveform_sig_loopback =7422;
25882: waveform_sig_loopback =7306;
25883: waveform_sig_loopback =6221;
25884: waveform_sig_loopback =8534;
25885: waveform_sig_loopback =6705;
25886: waveform_sig_loopback =6942;
25887: waveform_sig_loopback =7501;
25888: waveform_sig_loopback =7152;
25889: waveform_sig_loopback =7034;
25890: waveform_sig_loopback =6972;
25891: waveform_sig_loopback =8176;
25892: waveform_sig_loopback =6099;
25893: waveform_sig_loopback =7348;
25894: waveform_sig_loopback =7746;
25895: waveform_sig_loopback =6853;
25896: waveform_sig_loopback =6473;
25897: waveform_sig_loopback =8221;
25898: waveform_sig_loopback =6837;
25899: waveform_sig_loopback =5959;
25900: waveform_sig_loopback =8526;
25901: waveform_sig_loopback =7184;
25902: waveform_sig_loopback =5701;
25903: waveform_sig_loopback =7549;
25904: waveform_sig_loopback =8181;
25905: waveform_sig_loopback =6620;
25906: waveform_sig_loopback =5640;
25907: waveform_sig_loopback =8640;
25908: waveform_sig_loopback =7206;
25909: waveform_sig_loopback =6246;
25910: waveform_sig_loopback =8836;
25911: waveform_sig_loopback =3453;
25912: waveform_sig_loopback =8186;
25913: waveform_sig_loopback =9130;
25914: waveform_sig_loopback =5720;
25915: waveform_sig_loopback =6193;
25916: waveform_sig_loopback =6563;
25917: waveform_sig_loopback =8129;
25918: waveform_sig_loopback =7614;
25919: waveform_sig_loopback =5400;
25920: waveform_sig_loopback =7291;
25921: waveform_sig_loopback =7038;
25922: waveform_sig_loopback =6812;
25923: waveform_sig_loopback =7068;
25924: waveform_sig_loopback =5956;
25925: waveform_sig_loopback =7904;
25926: waveform_sig_loopback =6344;
25927: waveform_sig_loopback =6607;
25928: waveform_sig_loopback =7007;
25929: waveform_sig_loopback =6750;
25930: waveform_sig_loopback =6541;
25931: waveform_sig_loopback =6475;
25932: waveform_sig_loopback =7850;
25933: waveform_sig_loopback =5397;
25934: waveform_sig_loopback =6843;
25935: waveform_sig_loopback =7575;
25936: waveform_sig_loopback =5806;
25937: waveform_sig_loopback =6317;
25938: waveform_sig_loopback =7714;
25939: waveform_sig_loopback =6051;
25940: waveform_sig_loopback =5826;
25941: waveform_sig_loopback =7412;
25942: waveform_sig_loopback =6867;
25943: waveform_sig_loopback =5372;
25944: waveform_sig_loopback =6464;
25945: waveform_sig_loopback =7836;
25946: waveform_sig_loopback =5669;
25947: waveform_sig_loopback =5201;
25948: waveform_sig_loopback =8183;
25949: waveform_sig_loopback =5877;
25950: waveform_sig_loopback =6071;
25951: waveform_sig_loopback =7958;
25952: waveform_sig_loopback =2528;
25953: waveform_sig_loopback =7791;
25954: waveform_sig_loopback =8129;
25955: waveform_sig_loopback =5080;
25956: waveform_sig_loopback =5391;
25957: waveform_sig_loopback =5731;
25958: waveform_sig_loopback =7457;
25959: waveform_sig_loopback =6905;
25960: waveform_sig_loopback =4368;
25961: waveform_sig_loopback =6550;
25962: waveform_sig_loopback =6356;
25963: waveform_sig_loopback =5864;
25964: waveform_sig_loopback =6303;
25965: waveform_sig_loopback =5014;
25966: waveform_sig_loopback =7070;
25967: waveform_sig_loopback =5664;
25968: waveform_sig_loopback =5491;
25969: waveform_sig_loopback =6120;
25970: waveform_sig_loopback =6126;
25971: waveform_sig_loopback =5284;
25972: waveform_sig_loopback =5914;
25973: waveform_sig_loopback =6834;
25974: waveform_sig_loopback =4239;
25975: waveform_sig_loopback =6407;
25976: waveform_sig_loopback =6184;
25977: waveform_sig_loopback =4977;
25978: waveform_sig_loopback =5539;
25979: waveform_sig_loopback =6416;
25980: waveform_sig_loopback =5300;
25981: waveform_sig_loopback =4681;
25982: waveform_sig_loopback =6350;
25983: waveform_sig_loopback =5976;
25984: waveform_sig_loopback =4057;
25985: waveform_sig_loopback =5545;
25986: waveform_sig_loopback =6883;
25987: waveform_sig_loopback =4260;
25988: waveform_sig_loopback =4371;
25989: waveform_sig_loopback =7121;
25990: waveform_sig_loopback =4458;
25991: waveform_sig_loopback =5432;
25992: waveform_sig_loopback =6417;
25993: waveform_sig_loopback =1392;
25994: waveform_sig_loopback =7085;
25995: waveform_sig_loopback =6596;
25996: waveform_sig_loopback =4059;
25997: waveform_sig_loopback =4286;
25998: waveform_sig_loopback =4425;
25999: waveform_sig_loopback =6563;
26000: waveform_sig_loopback =5579;
26001: waveform_sig_loopback =3029;
26002: waveform_sig_loopback =5750;
26003: waveform_sig_loopback =4813;
26004: waveform_sig_loopback =4822;
26005: waveform_sig_loopback =5156;
26006: waveform_sig_loopback =3477;
26007: waveform_sig_loopback =6197;
26008: waveform_sig_loopback =4186;
26009: waveform_sig_loopback =4151;
26010: waveform_sig_loopback =5120;
26011: waveform_sig_loopback =4559;
26012: waveform_sig_loopback =4003;
26013: waveform_sig_loopback =4810;
26014: waveform_sig_loopback =5113;
26015: waveform_sig_loopback =3128;
26016: waveform_sig_loopback =5057;
26017: waveform_sig_loopback =4586;
26018: waveform_sig_loopback =3885;
26019: waveform_sig_loopback =3928;
26020: waveform_sig_loopback =5081;
26021: waveform_sig_loopback =4005;
26022: waveform_sig_loopback =3052;
26023: waveform_sig_loopback =5212;
26024: waveform_sig_loopback =4453;
26025: waveform_sig_loopback =2487;
26026: waveform_sig_loopback =4498;
26027: waveform_sig_loopback =5247;
26028: waveform_sig_loopback =2742;
26029: waveform_sig_loopback =3223;
26030: waveform_sig_loopback =5456;
26031: waveform_sig_loopback =3030;
26032: waveform_sig_loopback =4237;
26033: waveform_sig_loopback =4581;
26034: waveform_sig_loopback =172;
26035: waveform_sig_loopback =5733;
26036: waveform_sig_loopback =4883;
26037: waveform_sig_loopback =2791;
26038: waveform_sig_loopback =2542;
26039: waveform_sig_loopback =3047;
26040: waveform_sig_loopback =5239;
26041: waveform_sig_loopback =3636;
26042: waveform_sig_loopback =1694;
26043: waveform_sig_loopback =4216;
26044: waveform_sig_loopback =3005;
26045: waveform_sig_loopback =3594;
26046: waveform_sig_loopback =3209;
26047: waveform_sig_loopback =2014;
26048: waveform_sig_loopback =4856;
26049: waveform_sig_loopback =2129;
26050: waveform_sig_loopback =2868;
26051: waveform_sig_loopback =3438;
26052: waveform_sig_loopback =2771;
26053: waveform_sig_loopback =2590;
26054: waveform_sig_loopback =3035;
26055: waveform_sig_loopback =3430;
26056: waveform_sig_loopback =1672;
26057: waveform_sig_loopback =3207;
26058: waveform_sig_loopback =3051;
26059: waveform_sig_loopback =2244;
26060: waveform_sig_loopback =2169;
26061: waveform_sig_loopback =3632;
26062: waveform_sig_loopback =2141;
26063: waveform_sig_loopback =1362;
26064: waveform_sig_loopback =3879;
26065: waveform_sig_loopback =2437;
26066: waveform_sig_loopback =893;
26067: waveform_sig_loopback =3049;
26068: waveform_sig_loopback =3195;
26069: waveform_sig_loopback =1252;
26070: waveform_sig_loopback =1478;
26071: waveform_sig_loopback =3678;
26072: waveform_sig_loopback =1423;
26073: waveform_sig_loopback =2409;
26074: waveform_sig_loopback =2722;
26075: waveform_sig_loopback =-1484;
26076: waveform_sig_loopback =4006;
26077: waveform_sig_loopback =3116;
26078: waveform_sig_loopback =896;
26079: waveform_sig_loopback =700;
26080: waveform_sig_loopback =1474;
26081: waveform_sig_loopback =3371;
26082: waveform_sig_loopback =1690;
26083: waveform_sig_loopback =99;
26084: waveform_sig_loopback =2352;
26085: waveform_sig_loopback =1132;
26086: waveform_sig_loopback =2016;
26087: waveform_sig_loopback =1073;
26088: waveform_sig_loopback =568;
26089: waveform_sig_loopback =2920;
26090: waveform_sig_loopback =112;
26091: waveform_sig_loopback =1484;
26092: waveform_sig_loopback =1256;
26093: waveform_sig_loopback =1102;
26094: waveform_sig_loopback =882;
26095: waveform_sig_loopback =982;
26096: waveform_sig_loopback =1859;
26097: waveform_sig_loopback =-347;
26098: waveform_sig_loopback =1428;
26099: waveform_sig_loopback =1456;
26100: waveform_sig_loopback =-2;
26101: waveform_sig_loopback =606;
26102: waveform_sig_loopback =1807;
26103: waveform_sig_loopback =11;
26104: waveform_sig_loopback =-165;
26105: waveform_sig_loopback =1818;
26106: waveform_sig_loopback =570;
26107: waveform_sig_loopback =-867;
26108: waveform_sig_loopback =1116;
26109: waveform_sig_loopback =1335;
26110: waveform_sig_loopback =-652;
26111: waveform_sig_loopback =-366;
26112: waveform_sig_loopback =1851;
26113: waveform_sig_loopback =-524;
26114: waveform_sig_loopback =547;
26115: waveform_sig_loopback =770;
26116: waveform_sig_loopback =-3300;
26117: waveform_sig_loopback =2137;
26118: waveform_sig_loopback =1311;
26119: waveform_sig_loopback =-1168;
26120: waveform_sig_loopback =-1182;
26121: waveform_sig_loopback =-123;
26122: waveform_sig_loopback =1188;
26123: waveform_sig_loopback =-22;
26124: waveform_sig_loopback =-1815;
26125: waveform_sig_loopback =277;
26126: waveform_sig_loopback =-398;
26127: waveform_sig_loopback =-180;
26128: waveform_sig_loopback =-799;
26129: waveform_sig_loopback =-1080;
26130: waveform_sig_loopback =642;
26131: waveform_sig_loopback =-1436;
26132: waveform_sig_loopback =-573;
26133: waveform_sig_loopback =-781;
26134: waveform_sig_loopback =-417;
26135: waveform_sig_loopback =-1441;
26136: waveform_sig_loopback =-625;
26137: waveform_sig_loopback =-85;
26138: waveform_sig_loopback =-2428;
26139: waveform_sig_loopback =-175;
26140: waveform_sig_loopback =-684;
26141: waveform_sig_loopback =-1892;
26142: waveform_sig_loopback =-1114;
26143: waveform_sig_loopback =-207;
26144: waveform_sig_loopback =-1923;
26145: waveform_sig_loopback =-1906;
26146: waveform_sig_loopback =-115;
26147: waveform_sig_loopback =-1475;
26148: waveform_sig_loopback =-2642;
26149: waveform_sig_loopback =-826;
26150: waveform_sig_loopback =-521;
26151: waveform_sig_loopback =-2557;
26152: waveform_sig_loopback =-2383;
26153: waveform_sig_loopback =233;
26154: waveform_sig_loopback =-2692;
26155: waveform_sig_loopback =-1178;
26156: waveform_sig_loopback =-1106;
26157: waveform_sig_loopback =-5408;
26158: waveform_sig_loopback =679;
26159: waveform_sig_loopback =-743;
26160: waveform_sig_loopback =-3322;
26161: waveform_sig_loopback =-2647;
26162: waveform_sig_loopback =-2199;
26163: waveform_sig_loopback =-686;
26164: waveform_sig_loopback =-1764;
26165: waveform_sig_loopback =-4011;
26166: waveform_sig_loopback =-1178;
26167: waveform_sig_loopback =-2455;
26168: waveform_sig_loopback =-2160;
26169: waveform_sig_loopback =-2340;
26170: waveform_sig_loopback =-3203;
26171: waveform_sig_loopback =-1132;
26172: waveform_sig_loopback =-3221;
26173: waveform_sig_loopback =-2634;
26174: waveform_sig_loopback =-2339;
26175: waveform_sig_loopback =-2492;
26176: waveform_sig_loopback =-3312;
26177: waveform_sig_loopback =-2179;
26178: waveform_sig_loopback =-2223;
26179: waveform_sig_loopback =-4127;
26180: waveform_sig_loopback =-1992;
26181: waveform_sig_loopback =-2563;
26182: waveform_sig_loopback =-3718;
26183: waveform_sig_loopback =-2853;
26184: waveform_sig_loopback =-2123;
26185: waveform_sig_loopback =-3837;
26186: waveform_sig_loopback =-3479;
26187: waveform_sig_loopback =-2144;
26188: waveform_sig_loopback =-3138;
26189: waveform_sig_loopback =-4458;
26190: waveform_sig_loopback =-2695;
26191: waveform_sig_loopback =-2015;
26192: waveform_sig_loopback =-4726;
26193: waveform_sig_loopback =-3850;
26194: waveform_sig_loopback =-1459;
26195: waveform_sig_loopback =-4955;
26196: waveform_sig_loopback =-2187;
26197: waveform_sig_loopback =-3445;
26198: waveform_sig_loopback =-7097;
26199: waveform_sig_loopback =-589;
26200: waveform_sig_loopback =-3183;
26201: waveform_sig_loopback =-4598;
26202: waveform_sig_loopback =-4555;
26203: waveform_sig_loopback =-4065;
26204: waveform_sig_loopback =-1949;
26205: waveform_sig_loopback =-4032;
26206: waveform_sig_loopback =-5426;
26207: waveform_sig_loopback =-2781;
26208: waveform_sig_loopback =-4435;
26209: waveform_sig_loopback =-3572;
26210: waveform_sig_loopback =-4278;
26211: waveform_sig_loopback =-4777;
26212: waveform_sig_loopback =-2699;
26213: waveform_sig_loopback =-5093;
26214: waveform_sig_loopback =-4194;
26215: waveform_sig_loopback =-3990;
26216: waveform_sig_loopback =-4073;
26217: waveform_sig_loopback =-5106;
26218: waveform_sig_loopback =-3611;
26219: waveform_sig_loopback =-4040;
26220: waveform_sig_loopback =-5707;
26221: waveform_sig_loopback =-3290;
26222: waveform_sig_loopback =-4658;
26223: waveform_sig_loopback =-4949;
26224: waveform_sig_loopback =-4503;
26225: waveform_sig_loopback =-3918;
26226: waveform_sig_loopback =-5016;
26227: waveform_sig_loopback =-5510;
26228: waveform_sig_loopback =-3296;
26229: waveform_sig_loopback =-4803;
26230: waveform_sig_loopback =-6268;
26231: waveform_sig_loopback =-3695;
26232: waveform_sig_loopback =-3988;
26233: waveform_sig_loopback =-6275;
26234: waveform_sig_loopback =-5061;
26235: waveform_sig_loopback =-3253;
26236: waveform_sig_loopback =-6287;
26237: waveform_sig_loopback =-3693;
26238: waveform_sig_loopback =-5337;
26239: waveform_sig_loopback =-8155;
26240: waveform_sig_loopback =-2131;
26241: waveform_sig_loopback =-4807;
26242: waveform_sig_loopback =-5896;
26243: waveform_sig_loopback =-6183;
26244: waveform_sig_loopback =-5331;
26245: waveform_sig_loopback =-3285;
26246: waveform_sig_loopback =-5829;
26247: waveform_sig_loopback =-6617;
26248: waveform_sig_loopback =-4231;
26249: waveform_sig_loopback =-6197;
26250: waveform_sig_loopback =-4570;
26251: waveform_sig_loopback =-5925;
26252: waveform_sig_loopback =-6071;
26253: waveform_sig_loopback =-4204;
26254: waveform_sig_loopback =-6582;
26255: waveform_sig_loopback =-5230;
26256: waveform_sig_loopback =-5470;
26257: waveform_sig_loopback =-5690;
26258: waveform_sig_loopback =-6317;
26259: waveform_sig_loopback =-4685;
26260: waveform_sig_loopback =-5810;
26261: waveform_sig_loopback =-6788;
26262: waveform_sig_loopback =-4860;
26263: waveform_sig_loopback =-5899;
26264: waveform_sig_loopback =-6075;
26265: waveform_sig_loopback =-6324;
26266: waveform_sig_loopback =-4681;
26267: waveform_sig_loopback =-6608;
26268: waveform_sig_loopback =-6831;
26269: waveform_sig_loopback =-4318;
26270: waveform_sig_loopback =-6562;
26271: waveform_sig_loopback =-7121;
26272: waveform_sig_loopback =-5001;
26273: waveform_sig_loopback =-5518;
26274: waveform_sig_loopback =-7234;
26275: waveform_sig_loopback =-6362;
26276: waveform_sig_loopback =-4505;
26277: waveform_sig_loopback =-7509;
26278: waveform_sig_loopback =-4819;
26279: waveform_sig_loopback =-6663;
26280: waveform_sig_loopback =-9162;
26281: waveform_sig_loopback =-3254;
26282: waveform_sig_loopback =-6031;
26283: waveform_sig_loopback =-7034;
26284: waveform_sig_loopback =-7485;
26285: waveform_sig_loopback =-6241;
26286: waveform_sig_loopback =-4383;
26287: waveform_sig_loopback =-7146;
26288: waveform_sig_loopback =-7382;
26289: waveform_sig_loopback =-5492;
26290: waveform_sig_loopback =-6988;
26291: waveform_sig_loopback =-5600;
26292: waveform_sig_loopback =-7405;
26293: waveform_sig_loopback =-6614;
26294: waveform_sig_loopback =-5216;
26295: waveform_sig_loopback =-7763;
26296: waveform_sig_loopback =-6066;
26297: waveform_sig_loopback =-6635;
26298: waveform_sig_loopback =-6523;
26299: waveform_sig_loopback =-7181;
26300: waveform_sig_loopback =-6044;
26301: waveform_sig_loopback =-6510;
26302: waveform_sig_loopback =-7667;
26303: waveform_sig_loopback =-5899;
26304: waveform_sig_loopback =-6585;
26305: waveform_sig_loopback =-7320;
26306: waveform_sig_loopback =-6853;
26307: waveform_sig_loopback =-5650;
26308: waveform_sig_loopback =-7809;
26309: waveform_sig_loopback =-7255;
26310: waveform_sig_loopback =-5240;
26311: waveform_sig_loopback =-7541;
26312: waveform_sig_loopback =-7845;
26313: waveform_sig_loopback =-5779;
26314: waveform_sig_loopback =-6366;
26315: waveform_sig_loopback =-8030;
26316: waveform_sig_loopback =-7137;
26317: waveform_sig_loopback =-5230;
26318: waveform_sig_loopback =-8172;
26319: waveform_sig_loopback =-5649;
26320: waveform_sig_loopback =-7561;
26321: waveform_sig_loopback =-9611;
26322: waveform_sig_loopback =-4142;
26323: waveform_sig_loopback =-6632;
26324: waveform_sig_loopback =-7891;
26325: waveform_sig_loopback =-8142;
26326: waveform_sig_loopback =-6558;
26327: waveform_sig_loopback =-5513;
26328: waveform_sig_loopback =-7625;
26329: waveform_sig_loopback =-8025;
26330: waveform_sig_loopback =-6348;
26331: waveform_sig_loopback =-7295;
26332: waveform_sig_loopback =-6500;
26333: waveform_sig_loopback =-7917;
26334: waveform_sig_loopback =-7038;
26335: waveform_sig_loopback =-6170;
26336: waveform_sig_loopback =-8106;
26337: waveform_sig_loopback =-6742;
26338: waveform_sig_loopback =-7255;
26339: waveform_sig_loopback =-6877;
26340: waveform_sig_loopback =-7827;
26341: waveform_sig_loopback =-6438;
26342: waveform_sig_loopback =-7065;
26343: waveform_sig_loopback =-8201;
26344: waveform_sig_loopback =-6331;
26345: waveform_sig_loopback =-6978;
26346: waveform_sig_loopback =-7972;
26347: waveform_sig_loopback =-7031;
26348: waveform_sig_loopback =-6146;
26349: waveform_sig_loopback =-8391;
26350: waveform_sig_loopback =-7291;
26351: waveform_sig_loopback =-5948;
26352: waveform_sig_loopback =-7908;
26353: waveform_sig_loopback =-8017;
26354: waveform_sig_loopback =-6352;
26355: waveform_sig_loopback =-6511;
26356: waveform_sig_loopback =-8462;
26357: waveform_sig_loopback =-7499;
26358: waveform_sig_loopback =-5359;
26359: waveform_sig_loopback =-8763;
26360: waveform_sig_loopback =-5711;
26361: waveform_sig_loopback =-7938;
26362: waveform_sig_loopback =-9989;
26363: waveform_sig_loopback =-4042;
26364: waveform_sig_loopback =-7097;
26365: waveform_sig_loopback =-8317;
26366: waveform_sig_loopback =-8027;
26367: waveform_sig_loopback =-6911;
26368: waveform_sig_loopback =-5696;
26369: waveform_sig_loopback =-7720;
26370: waveform_sig_loopback =-8349;
26371: waveform_sig_loopback =-6292;
26372: waveform_sig_loopback =-7515;
26373: waveform_sig_loopback =-6813;
26374: waveform_sig_loopback =-7772;
26375: waveform_sig_loopback =-7255;
26376: waveform_sig_loopback =-6340;
26377: waveform_sig_loopback =-8008;
26378: waveform_sig_loopback =-6966;
26379: waveform_sig_loopback =-7212;
26380: waveform_sig_loopback =-6922;
26381: waveform_sig_loopback =-8059;
26382: waveform_sig_loopback =-6237;
26383: waveform_sig_loopback =-7174;
26384: waveform_sig_loopback =-8273;
26385: waveform_sig_loopback =-6085;
26386: waveform_sig_loopback =-7215;
26387: waveform_sig_loopback =-7956;
26388: waveform_sig_loopback =-6684;
26389: waveform_sig_loopback =-6457;
26390: waveform_sig_loopback =-8193;
26391: waveform_sig_loopback =-7079;
26392: waveform_sig_loopback =-6103;
26393: waveform_sig_loopback =-7535;
26394: waveform_sig_loopback =-8092;
26395: waveform_sig_loopback =-6133;
26396: waveform_sig_loopback =-6266;
26397: waveform_sig_loopback =-8698;
26398: waveform_sig_loopback =-6888;
26399: waveform_sig_loopback =-5348;
26400: waveform_sig_loopback =-8774;
26401: waveform_sig_loopback =-5080;
26402: waveform_sig_loopback =-8248;
26403: waveform_sig_loopback =-9491;
26404: waveform_sig_loopback =-3690;
26405: waveform_sig_loopback =-7165;
26406: waveform_sig_loopback =-7875;
26407: waveform_sig_loopback =-7745;
26408: waveform_sig_loopback =-6734;
26409: waveform_sig_loopback =-5183;
26410: waveform_sig_loopback =-7641;
26411: waveform_sig_loopback =-8036;
26412: waveform_sig_loopback =-5755;
26413: waveform_sig_loopback =-7399;
26414: waveform_sig_loopback =-6345;
26415: waveform_sig_loopback =-7435;
26416: waveform_sig_loopback =-6979;
26417: waveform_sig_loopback =-5823;
26418: waveform_sig_loopback =-7640;
26419: waveform_sig_loopback =-6672;
26420: waveform_sig_loopback =-6586;
26421: waveform_sig_loopback =-6594;
26422: waveform_sig_loopback =-7653;
26423: waveform_sig_loopback =-5451;
26424: waveform_sig_loopback =-7161;
26425: waveform_sig_loopback =-7511;
26426: waveform_sig_loopback =-5484;
26427: waveform_sig_loopback =-7061;
26428: waveform_sig_loopback =-6981;
26429: waveform_sig_loopback =-6400;
26430: waveform_sig_loopback =-5907;
26431: waveform_sig_loopback =-7437;
26432: waveform_sig_loopback =-6770;
26433: waveform_sig_loopback =-5272;
26434: waveform_sig_loopback =-7130;
26435: waveform_sig_loopback =-7561;
26436: waveform_sig_loopback =-5215;
26437: waveform_sig_loopback =-5909;
26438: waveform_sig_loopback =-8104;
26439: waveform_sig_loopback =-5957;
26440: waveform_sig_loopback =-4972;
26441: waveform_sig_loopback =-8043;
26442: waveform_sig_loopback =-4185;
26443: waveform_sig_loopback =-8014;
26444: waveform_sig_loopback =-8365;
26445: waveform_sig_loopback =-2982;
26446: waveform_sig_loopback =-6712;
26447: waveform_sig_loopback =-6880;
26448: waveform_sig_loopback =-7205;
26449: waveform_sig_loopback =-5896;
26450: waveform_sig_loopback =-4197;
26451: waveform_sig_loopback =-7283;
26452: waveform_sig_loopback =-7011;
26453: waveform_sig_loopback =-4934;
26454: waveform_sig_loopback =-6883;
26455: waveform_sig_loopback =-5121;
26456: waveform_sig_loopback =-6977;
26457: waveform_sig_loopback =-6009;
26458: waveform_sig_loopback =-4790;
26459: waveform_sig_loopback =-7157;
26460: waveform_sig_loopback =-5519;
26461: waveform_sig_loopback =-5747;
26462: waveform_sig_loopback =-5944;
26463: waveform_sig_loopback =-6435;
26464: waveform_sig_loopback =-4696;
26465: waveform_sig_loopback =-6364;
26466: waveform_sig_loopback =-6250;
26467: waveform_sig_loopback =-4803;
26468: waveform_sig_loopback =-5994;
26469: waveform_sig_loopback =-5988;
26470: waveform_sig_loopback =-5547;
26471: waveform_sig_loopback =-4725;
26472: waveform_sig_loopback =-6555;
26473: waveform_sig_loopback =-5788;
26474: waveform_sig_loopback =-4043;
26475: waveform_sig_loopback =-6291;
26476: waveform_sig_loopback =-6466;
26477: waveform_sig_loopback =-3968;
26478: waveform_sig_loopback =-5181;
26479: waveform_sig_loopback =-6850;
26480: waveform_sig_loopback =-4729;
26481: waveform_sig_loopback =-4243;
26482: waveform_sig_loopback =-6568;
26483: waveform_sig_loopback =-3202;
26484: waveform_sig_loopback =-7185;
26485: waveform_sig_loopback =-6682;
26486: waveform_sig_loopback =-2207;
26487: waveform_sig_loopback =-5397;
26488: waveform_sig_loopback =-5700;
26489: waveform_sig_loopback =-6278;
26490: waveform_sig_loopback =-4247;
26491: waveform_sig_loopback =-3218;
26492: waveform_sig_loopback =-6194;
26493: waveform_sig_loopback =-5432;
26494: waveform_sig_loopback =-3978;
26495: waveform_sig_loopback =-5442;
26496: waveform_sig_loopback =-3793;
26497: waveform_sig_loopback =-6016;
26498: waveform_sig_loopback =-4320;
26499: waveform_sig_loopback =-3670;
26500: waveform_sig_loopback =-5971;
26501: waveform_sig_loopback =-3915;
26502: waveform_sig_loopback =-4673;
26503: waveform_sig_loopback =-4566;
26504: waveform_sig_loopback =-4927;
26505: waveform_sig_loopback =-3620;
26506: waveform_sig_loopback =-4810;
26507: waveform_sig_loopback =-4901;
26508: waveform_sig_loopback =-3656;
26509: waveform_sig_loopback =-4358;
26510: waveform_sig_loopback =-4851;
26511: waveform_sig_loopback =-4021;
26512: waveform_sig_loopback =-3271;
26513: waveform_sig_loopback =-5477;
26514: waveform_sig_loopback =-4060;
26515: waveform_sig_loopback =-2676;
26516: waveform_sig_loopback =-5161;
26517: waveform_sig_loopback =-4715;
26518: waveform_sig_loopback =-2619;
26519: waveform_sig_loopback =-3899;
26520: waveform_sig_loopback =-5185;
26521: waveform_sig_loopback =-3410;
26522: waveform_sig_loopback =-2728;
26523: waveform_sig_loopback =-4964;
26524: waveform_sig_loopback =-1971;
26525: waveform_sig_loopback =-5648;
26526: waveform_sig_loopback =-5061;
26527: waveform_sig_loopback =-811;
26528: waveform_sig_loopback =-3730;
26529: waveform_sig_loopback =-4508;
26530: waveform_sig_loopback =-4560;
26531: waveform_sig_loopback =-2574;
26532: waveform_sig_loopback =-2054;
26533: waveform_sig_loopback =-4447;
26534: waveform_sig_loopback =-3882;
26535: waveform_sig_loopback =-2625;
26536: waveform_sig_loopback =-3644;
26537: waveform_sig_loopback =-2382;
26538: waveform_sig_loopback =-4428;
26539: waveform_sig_loopback =-2515;
26540: waveform_sig_loopback =-2468;
26541: waveform_sig_loopback =-4174;
26542: waveform_sig_loopback =-2167;
26543: waveform_sig_loopback =-3364;
26544: waveform_sig_loopback =-2729;
26545: waveform_sig_loopback =-3413;
26546: waveform_sig_loopback =-1951;
26547: waveform_sig_loopback =-2969;
26548: waveform_sig_loopback =-3653;
26549: waveform_sig_loopback =-1728;
26550: waveform_sig_loopback =-2550;
26551: waveform_sig_loopback =-3509;
26552: waveform_sig_loopback =-2002;
26553: waveform_sig_loopback =-1893;
26554: waveform_sig_loopback =-3732;
26555: waveform_sig_loopback =-1979;
26556: waveform_sig_loopback =-1409;
26557: waveform_sig_loopback =-3277;
26558: waveform_sig_loopback =-2963;
26559: waveform_sig_loopback =-1028;
26560: waveform_sig_loopback =-2015;
26561: waveform_sig_loopback =-3614;
26562: waveform_sig_loopback =-1547;
26563: waveform_sig_loopback =-1011;
26564: waveform_sig_loopback =-3278;
26565: waveform_sig_loopback =-83;
26566: waveform_sig_loopback =-3997;
26567: waveform_sig_loopback =-3262;
26568: waveform_sig_loopback =1032;
26569: waveform_sig_loopback =-1913;
26570: waveform_sig_loopback =-2968;
26571: waveform_sig_loopback =-2517;
26572: waveform_sig_loopback =-851;
26573: waveform_sig_loopback =-354;
26574: waveform_sig_loopback =-2462;
26575: waveform_sig_loopback =-2306;
26576: waveform_sig_loopback =-652;
26577: waveform_sig_loopback =-1717;
26578: waveform_sig_loopback =-934;
26579: waveform_sig_loopback =-2281;
26580: waveform_sig_loopback =-743;
26581: waveform_sig_loopback =-835;
26582: waveform_sig_loopback =-2009;
26583: waveform_sig_loopback =-805;
26584: waveform_sig_loopback =-1200;
26585: waveform_sig_loopback =-858;
26586: waveform_sig_loopback =-1913;
26587: waveform_sig_loopback =291;
26588: waveform_sig_loopback =-1568;
26589: waveform_sig_loopback =-1508;
26590: waveform_sig_loopback =293;
26591: waveform_sig_loopback =-1164;
26592: waveform_sig_loopback =-1367;
26593: waveform_sig_loopback =-129;
26594: waveform_sig_loopback =-194;
26595: waveform_sig_loopback =-1782;
26596: waveform_sig_loopback =-247;
26597: waveform_sig_loopback =419;
26598: waveform_sig_loopback =-1613;
26599: waveform_sig_loopback =-905;
26600: waveform_sig_loopback =879;
26601: waveform_sig_loopback =-282;
26602: waveform_sig_loopback =-1996;
26603: waveform_sig_loopback =577;
26604: waveform_sig_loopback =1077;
26605: waveform_sig_loopback =-1806;
26606: waveform_sig_loopback =1921;
26607: waveform_sig_loopback =-2363;
26608: waveform_sig_loopback =-1098;
26609: waveform_sig_loopback =3132;
26610: waveform_sig_loopback =-682;
26611: waveform_sig_loopback =-822;
26612: waveform_sig_loopback =-386;
26613: waveform_sig_loopback =645;
26614: waveform_sig_loopback =1837;
26615: waveform_sig_loopback =-875;
26616: waveform_sig_loopback =-302;
26617: waveform_sig_loopback =1401;
26618: waveform_sig_loopback =-304;
26619: waveform_sig_loopback =1321;
26620: waveform_sig_loopback =-455;
26621: waveform_sig_loopback =897;
26622: waveform_sig_loopback =1327;
26623: waveform_sig_loopback =-297;
26624: waveform_sig_loopback =1153;
26625: waveform_sig_loopback =775;
26626: waveform_sig_loopback =673;
26627: waveform_sig_loopback =353;
26628: waveform_sig_loopback =2109;
26629: waveform_sig_loopback =97;
26630: waveform_sig_loopback =577;
26631: waveform_sig_loopback =2039;
26632: waveform_sig_loopback =701;
26633: waveform_sig_loopback =490;
26634: waveform_sig_loopback =1834;
26635: waveform_sig_loopback =1606;
26636: waveform_sig_loopback =180;
26637: waveform_sig_loopback =1623;
26638: waveform_sig_loopback =2281;
26639: waveform_sig_loopback =593;
26640: waveform_sig_loopback =647;
26641: waveform_sig_loopback =2915;
26642: waveform_sig_loopback =1627;
26643: waveform_sig_loopback =-136;
26644: waveform_sig_loopback =2794;
26645: waveform_sig_loopback =2353;
26646: waveform_sig_loopback =343;
26647: waveform_sig_loopback =4218;
26648: waveform_sig_loopback =-1227;
26649: waveform_sig_loopback =1328;
26650: waveform_sig_loopback =4865;
26651: waveform_sig_loopback =970;
26652: waveform_sig_loopback =1504;
26653: waveform_sig_loopback =940;
26654: waveform_sig_loopback =2978;
26655: waveform_sig_loopback =3764;
26656: waveform_sig_loopback =444;
26657: waveform_sig_loopback =2153;
26658: waveform_sig_loopback =2902;
26659: waveform_sig_loopback =1735;
26660: waveform_sig_loopback =3249;
26661: waveform_sig_loopback =998;
26662: waveform_sig_loopback =3257;
26663: waveform_sig_loopback =2878;
26664: waveform_sig_loopback =1490;
26665: waveform_sig_loopback =3085;
26666: waveform_sig_loopback =2543;
26667: waveform_sig_loopback =2597;
26668: waveform_sig_loopback =2023;
26669: waveform_sig_loopback =4055;
26670: waveform_sig_loopback =1761;
26671: waveform_sig_loopback =2572;
26672: waveform_sig_loopback =3780;
26673: waveform_sig_loopback =2293;
26674: waveform_sig_loopback =2691;
26675: waveform_sig_loopback =3335;
26676: waveform_sig_loopback =3478;
26677: waveform_sig_loopback =2062;
26678: waveform_sig_loopback =3185;
26679: waveform_sig_loopback =4491;
26680: waveform_sig_loopback =1899;
26681: waveform_sig_loopback =2646;
26682: waveform_sig_loopback =4988;
26683: waveform_sig_loopback =2782;
26684: waveform_sig_loopback =2094;
26685: waveform_sig_loopback =4457;
26686: waveform_sig_loopback =3831;
26687: waveform_sig_loopback =2604;
26688: waveform_sig_loopback =5441;
26689: waveform_sig_loopback =646;
26690: waveform_sig_loopback =3388;
26691: waveform_sig_loopback =6193;
26692: waveform_sig_loopback =3095;
26693: waveform_sig_loopback =2912;
26694: waveform_sig_loopback =2703;
26695: waveform_sig_loopback =5021;
26696: waveform_sig_loopback =5096;
26697: waveform_sig_loopback =2288;
26698: waveform_sig_loopback =3885;
26699: waveform_sig_loopback =4417;
26700: waveform_sig_loopback =3654;
26701: waveform_sig_loopback =4758;
26702: waveform_sig_loopback =2597;
26703: waveform_sig_loopback =5117;
26704: waveform_sig_loopback =4371;
26705: waveform_sig_loopback =3228;
26706: waveform_sig_loopback =4748;
26707: waveform_sig_loopback =4151;
26708: waveform_sig_loopback =4136;
26709: waveform_sig_loopback =3931;
26710: waveform_sig_loopback =5402;
26711: waveform_sig_loopback =3317;
26712: waveform_sig_loopback =4523;
26713: waveform_sig_loopback =4967;
26714: waveform_sig_loopback =4316;
26715: waveform_sig_loopback =3875;
26716: waveform_sig_loopback =4988;
26717: waveform_sig_loopback =5402;
26718: waveform_sig_loopback =2983;
26719: waveform_sig_loopback =5364;
26720: waveform_sig_loopback =5817;
26721: waveform_sig_loopback =3226;
26722: waveform_sig_loopback =4713;
26723: waveform_sig_loopback =6085;
26724: waveform_sig_loopback =4551;
26725: waveform_sig_loopback =3699;
26726: waveform_sig_loopback =5785;
26727: waveform_sig_loopback =5575;
26728: waveform_sig_loopback =3994;
26729: waveform_sig_loopback =6962;
26730: waveform_sig_loopback =2121;
26731: waveform_sig_loopback =4940;
26732: waveform_sig_loopback =7767;
26733: waveform_sig_loopback =4437;
26734: waveform_sig_loopback =4235;
26735: waveform_sig_loopback =4387;
26736: waveform_sig_loopback =6454;
26737: waveform_sig_loopback =6410;
26738: waveform_sig_loopback =3733;
26739: waveform_sig_loopback =5458;
26740: waveform_sig_loopback =5670;
26741: waveform_sig_loopback =5198;
26742: waveform_sig_loopback =6077;
26743: waveform_sig_loopback =4029;
26744: waveform_sig_loopback =6745;
26745: waveform_sig_loopback =5442;
26746: waveform_sig_loopback =4796;
26747: waveform_sig_loopback =6314;
26748: waveform_sig_loopback =5245;
26749: waveform_sig_loopback =5700;
26750: waveform_sig_loopback =5195;
26751: waveform_sig_loopback =6718;
26752: waveform_sig_loopback =4971;
26753: waveform_sig_loopback =5454;
26754: waveform_sig_loopback =6604;
26755: waveform_sig_loopback =5574;
26756: waveform_sig_loopback =5006;
26757: waveform_sig_loopback =6740;
26758: waveform_sig_loopback =6169;
26759: waveform_sig_loopback =4517;
26760: waveform_sig_loopback =6860;
26761: waveform_sig_loopback =6607;
26762: waveform_sig_loopback =4752;
26763: waveform_sig_loopback =5951;
26764: waveform_sig_loopback =7209;
26765: waveform_sig_loopback =5843;
26766: waveform_sig_loopback =4705;
26767: waveform_sig_loopback =7282;
26768: waveform_sig_loopback =6600;
26769: waveform_sig_loopback =5120;
26770: waveform_sig_loopback =8219;
26771: waveform_sig_loopback =3091;
26772: waveform_sig_loopback =6378;
26773: waveform_sig_loopback =8727;
26774: waveform_sig_loopback =5552;
26775: waveform_sig_loopback =5331;
26776: waveform_sig_loopback =5608;
26777: waveform_sig_loopback =7591;
26778: waveform_sig_loopback =7237;
26779: waveform_sig_loopback =5078;
26780: waveform_sig_loopback =6378;
26781: waveform_sig_loopback =6777;
26782: waveform_sig_loopback =6443;
26783: waveform_sig_loopback =6740;
26784: waveform_sig_loopback =5468;
26785: waveform_sig_loopback =7632;
26786: waveform_sig_loopback =6305;
26787: waveform_sig_loopback =6170;
26788: waveform_sig_loopback =6808;
26789: waveform_sig_loopback =6568;
26790: waveform_sig_loopback =6648;
26791: waveform_sig_loopback =5937;
26792: waveform_sig_loopback =8058;
26793: waveform_sig_loopback =5460;
26794: waveform_sig_loopback =6636;
26795: waveform_sig_loopback =7626;
26796: waveform_sig_loopback =6160;
26797: waveform_sig_loopback =6239;
26798: waveform_sig_loopback =7596;
26799: waveform_sig_loopback =6935;
26800: waveform_sig_loopback =5511;
26801: waveform_sig_loopback =7682;
26802: waveform_sig_loopback =7407;
26803: waveform_sig_loopback =5634;
26804: waveform_sig_loopback =6781;
26805: waveform_sig_loopback =7992;
26806: waveform_sig_loopback =6711;
26807: waveform_sig_loopback =5376;
26808: waveform_sig_loopback =8247;
26809: waveform_sig_loopback =7307;
26810: waveform_sig_loopback =5817;
26811: waveform_sig_loopback =9163;
26812: waveform_sig_loopback =3525;
26813: waveform_sig_loopback =7328;
26814: waveform_sig_loopback =9570;
26815: waveform_sig_loopback =5887;
26816: waveform_sig_loopback =6192;
26817: waveform_sig_loopback =6423;
26818: waveform_sig_loopback =8113;
26819: waveform_sig_loopback =8109;
26820: waveform_sig_loopback =5529;
26821: waveform_sig_loopback =7072;
26822: waveform_sig_loopback =7600;
26823: waveform_sig_loopback =6803;
26824: waveform_sig_loopback =7451;
26825: waveform_sig_loopback =6157;
26826: waveform_sig_loopback =7986;
26827: waveform_sig_loopback =7080;
26828: waveform_sig_loopback =6655;
26829: waveform_sig_loopback =7279;
26830: waveform_sig_loopback =7417;
26831: waveform_sig_loopback =6829;
26832: waveform_sig_loopback =6728;
26833: waveform_sig_loopback =8571;
26834: waveform_sig_loopback =5705;
26835: waveform_sig_loopback =7460;
26836: waveform_sig_loopback =7952;
26837: waveform_sig_loopback =6531;
26838: waveform_sig_loopback =6883;
26839: waveform_sig_loopback =7894;
26840: waveform_sig_loopback =7316;
26841: waveform_sig_loopback =6074;
26842: waveform_sig_loopback =7943;
26843: waveform_sig_loopback =7857;
26844: waveform_sig_loopback =5969;
26845: waveform_sig_loopback =7074;
26846: waveform_sig_loopback =8506;
26847: waveform_sig_loopback =6871;
26848: waveform_sig_loopback =5679;
26849: waveform_sig_loopback =8844;
26850: waveform_sig_loopback =7246;
26851: waveform_sig_loopback =6332;
26852: waveform_sig_loopback =9462;
26853: waveform_sig_loopback =3415;
26854: waveform_sig_loopback =8107;
26855: waveform_sig_loopback =9636;
26856: waveform_sig_loopback =5958;
26857: waveform_sig_loopback =6693;
26858: waveform_sig_loopback =6422;
26859: waveform_sig_loopback =8470;
26860: waveform_sig_loopback =8346;
26861: waveform_sig_loopback =5373;
26862: waveform_sig_loopback =7633;
26863: waveform_sig_loopback =7611;
26864: waveform_sig_loopback =6860;
26865: waveform_sig_loopback =7802;
26866: waveform_sig_loopback =6012;
26867: waveform_sig_loopback =8261;
26868: waveform_sig_loopback =7207;
26869: waveform_sig_loopback =6472;
26870: waveform_sig_loopback =7588;
26871: waveform_sig_loopback =7386;
26872: waveform_sig_loopback =6707;
26873: waveform_sig_loopback =7049;
26874: waveform_sig_loopback =8344;
26875: waveform_sig_loopback =5747;
26876: waveform_sig_loopback =7645;
26877: waveform_sig_loopback =7638;
26878: waveform_sig_loopback =6663;
26879: waveform_sig_loopback =6899;
26880: waveform_sig_loopback =7718;
26881: waveform_sig_loopback =7325;
26882: waveform_sig_loopback =5898;
26883: waveform_sig_loopback =7927;
26884: waveform_sig_loopback =7855;
26885: waveform_sig_loopback =5583;
26886: waveform_sig_loopback =7129;
26887: waveform_sig_loopback =8538;
26888: waveform_sig_loopback =6384;
26889: waveform_sig_loopback =5730;
26890: waveform_sig_loopback =8706;
26891: waveform_sig_loopback =6806;
26892: waveform_sig_loopback =6608;
26893: waveform_sig_loopback =8825;
26894: waveform_sig_loopback =3252;
26895: waveform_sig_loopback =8306;
26896: waveform_sig_loopback =8979;
26897: waveform_sig_loopback =5875;
26898: waveform_sig_loopback =6433;
26899: waveform_sig_loopback =6108;
26900: waveform_sig_loopback =8437;
26901: waveform_sig_loopback =7805;
26902: waveform_sig_loopback =5027;
26903: waveform_sig_loopback =7719;
26904: waveform_sig_loopback =6880;
26905: waveform_sig_loopback =6718;
26906: waveform_sig_loopback =7508;
26907: waveform_sig_loopback =5487;
26908: waveform_sig_loopback =8216;
26909: waveform_sig_loopback =6481;
26910: waveform_sig_loopback =6221;
26911: waveform_sig_loopback =7384;
26912: waveform_sig_loopback =6644;
26913: waveform_sig_loopback =6454;
26914: waveform_sig_loopback =6747;
26915: waveform_sig_loopback =7604;
26916: waveform_sig_loopback =5393;
26917: waveform_sig_loopback =7234;
26918: waveform_sig_loopback =7135;
26919: waveform_sig_loopback =6099;
26920: waveform_sig_loopback =6290;
26921: waveform_sig_loopback =7393;
26922: waveform_sig_loopback =6704;
26923: waveform_sig_loopback =5316;
26924: waveform_sig_loopback =7447;
26925: waveform_sig_loopback =7343;
26926: waveform_sig_loopback =4920;
26927: waveform_sig_loopback =6655;
26928: waveform_sig_loopback =7985;
26929: waveform_sig_loopback =5458;
26930: waveform_sig_loopback =5525;
26931: waveform_sig_loopback =7978;
26932: waveform_sig_loopback =5930;
26933: waveform_sig_loopback =6360;
26934: waveform_sig_loopback =7724;
26935: waveform_sig_loopback =2792;
26936: waveform_sig_loopback =7742;
26937: waveform_sig_loopback =7873;
26938: waveform_sig_loopback =5632;
26939: waveform_sig_loopback =5205;
26940: waveform_sig_loopback =5450;
26941: waveform_sig_loopback =8003;
26942: waveform_sig_loopback =6664;
26943: waveform_sig_loopback =4441;
26944: waveform_sig_loopback =6735;
26945: waveform_sig_loopback =6067;
26946: waveform_sig_loopback =6246;
26947: waveform_sig_loopback =6097;
26948: waveform_sig_loopback =4667;
26949: waveform_sig_loopback =7762;
26950: waveform_sig_loopback =5323;
26951: waveform_sig_loopback =5366;
26952: waveform_sig_loopback =6259;
26953: waveform_sig_loopback =5910;
26954: waveform_sig_loopback =5611;
26955: waveform_sig_loopback =5700;
26956: waveform_sig_loopback =6472;
26957: waveform_sig_loopback =4673;
26958: waveform_sig_loopback =6312;
26959: waveform_sig_loopback =5886;
26960: waveform_sig_loopback =5376;
26961: waveform_sig_loopback =5085;
26962: waveform_sig_loopback =6644;
26963: waveform_sig_loopback =5520;
26964: waveform_sig_loopback =4001;
26965: waveform_sig_loopback =7047;
26966: waveform_sig_loopback =5791;
26967: waveform_sig_loopback =3816;
26968: waveform_sig_loopback =5939;
26969: waveform_sig_loopback =6564;
26970: waveform_sig_loopback =4597;
26971: waveform_sig_loopback =4311;
26972: waveform_sig_loopback =6785;
26973: waveform_sig_loopback =5086;
26974: waveform_sig_loopback =5024;
26975: waveform_sig_loopback =6487;
26976: waveform_sig_loopback =1852;
26977: waveform_sig_loopback =6534;
26978: waveform_sig_loopback =6838;
26979: waveform_sig_loopback =4296;
26980: waveform_sig_loopback =3923;
26981: waveform_sig_loopback =4681;
26982: waveform_sig_loopback =6458;
26983: waveform_sig_loopback =5407;
26984: waveform_sig_loopback =3466;
26985: waveform_sig_loopback =5354;
26986: waveform_sig_loopback =4886;
26987: waveform_sig_loopback =4982;
26988: waveform_sig_loopback =4813;
26989: waveform_sig_loopback =3784;
26990: waveform_sig_loopback =6123;
26991: waveform_sig_loopback =3953;
26992: waveform_sig_loopback =4491;
26993: waveform_sig_loopback =4990;
26994: waveform_sig_loopback =4388;
26995: waveform_sig_loopback =4364;
26996: waveform_sig_loopback =4446;
26997: waveform_sig_loopback =5265;
26998: waveform_sig_loopback =3321;
26999: waveform_sig_loopback =4632;
27000: waveform_sig_loopback =5055;
27001: waveform_sig_loopback =3759;
27002: waveform_sig_loopback =3695;
27003: waveform_sig_loopback =5599;
27004: waveform_sig_loopback =3650;
27005: waveform_sig_loopback =3118;
27006: waveform_sig_loopback =5523;
27007: waveform_sig_loopback =4083;
27008: waveform_sig_loopback =2858;
27009: waveform_sig_loopback =4382;
27010: waveform_sig_loopback =5065;
27011: waveform_sig_loopback =3274;
27012: waveform_sig_loopback =2683;
27013: waveform_sig_loopback =5649;
27014: waveform_sig_loopback =3331;
27015: waveform_sig_loopback =3573;
27016: waveform_sig_loopback =5164;
27017: waveform_sig_loopback =79;
27018: waveform_sig_loopback =5310;
27019: waveform_sig_loopback =5285;
27020: waveform_sig_loopback =2607;
27021: waveform_sig_loopback =2549;
27022: waveform_sig_loopback =3223;
27023: waveform_sig_loopback =4873;
27024: waveform_sig_loopback =3877;
27025: waveform_sig_loopback =1898;
27026: waveform_sig_loopback =3729;
27027: waveform_sig_loopback =3470;
27028: waveform_sig_loopback =3357;
27029: waveform_sig_loopback =3119;
27030: waveform_sig_loopback =2493;
27031: waveform_sig_loopback =4278;
27032: waveform_sig_loopback =2454;
27033: waveform_sig_loopback =2999;
27034: waveform_sig_loopback =3063;
27035: waveform_sig_loopback =3176;
27036: waveform_sig_loopback =2488;
27037: waveform_sig_loopback =2811;
27038: waveform_sig_loopback =3920;
27039: waveform_sig_loopback =1280;
27040: waveform_sig_loopback =3342;
27041: waveform_sig_loopback =3365;
27042: waveform_sig_loopback =1766;
27043: waveform_sig_loopback =2510;
27044: waveform_sig_loopback =3588;
27045: waveform_sig_loopback =1938;
27046: waveform_sig_loopback =1739;
27047: waveform_sig_loopback =3470;
27048: waveform_sig_loopback =2611;
27049: waveform_sig_loopback =1023;
27050: waveform_sig_loopback =2621;
27051: waveform_sig_loopback =3554;
27052: waveform_sig_loopback =1258;
27053: waveform_sig_loopback =1117;
27054: waveform_sig_loopback =3984;
27055: waveform_sig_loopback =1461;
27056: waveform_sig_loopback =2004;
27057: waveform_sig_loopback =3297;
27058: waveform_sig_loopback =-1740;
27059: waveform_sig_loopback =3788;
27060: waveform_sig_loopback =3548;
27061: waveform_sig_loopback =519;
27062: waveform_sig_loopback =1045;
27063: waveform_sig_loopback =1370;
27064: waveform_sig_loopback =2967;
27065: waveform_sig_loopback =2398;
27066: waveform_sig_loopback =-327;
27067: waveform_sig_loopback =2254;
27068: waveform_sig_loopback =1680;
27069: waveform_sig_loopback =1305;
27070: waveform_sig_loopback =1630;
27071: waveform_sig_loopback =409;
27072: waveform_sig_loopback =2538;
27073: waveform_sig_loopback =801;
27074: waveform_sig_loopback =908;
27075: waveform_sig_loopback =1500;
27076: waveform_sig_loopback =1301;
27077: waveform_sig_loopback =440;
27078: waveform_sig_loopback =1386;
27079: waveform_sig_loopback =1764;
27080: waveform_sig_loopback =-513;
27081: waveform_sig_loopback =1695;
27082: waveform_sig_loopback =1266;
27083: waveform_sig_loopback =8;
27084: waveform_sig_loopback =727;
27085: waveform_sig_loopback =1611;
27086: waveform_sig_loopback =89;
27087: waveform_sig_loopback =-42;
27088: waveform_sig_loopback =1535;
27089: waveform_sig_loopback =858;
27090: waveform_sig_loopback =-918;
27091: waveform_sig_loopback =783;
27092: waveform_sig_loopback =1931;
27093: waveform_sig_loopback =-961;
27094: waveform_sig_loopback =-489;
27095: waveform_sig_loopback =2239;
27096: waveform_sig_loopback =-869;
27097: waveform_sig_loopback =658;
27098: waveform_sig_loopback =1000;
27099: waveform_sig_loopback =-3643;
27100: waveform_sig_loopback =2387;
27101: waveform_sig_loopback =1122;
27102: waveform_sig_loopback =-1116;
27103: waveform_sig_loopback =-764;
27104: waveform_sig_loopback =-780;
27105: waveform_sig_loopback =1540;
27106: waveform_sig_loopback =179;
27107: waveform_sig_loopback =-2268;
27108: waveform_sig_loopback =785;
27109: waveform_sig_loopback =-725;
27110: waveform_sig_loopback =-230;
27111: waveform_sig_loopback =-323;
27112: waveform_sig_loopback =-1697;
27113: waveform_sig_loopback =1021;
27114: waveform_sig_loopback =-1451;
27115: waveform_sig_loopback =-856;
27116: waveform_sig_loopback =-297;
27117: waveform_sig_loopback =-800;
27118: waveform_sig_loopback =-1317;
27119: waveform_sig_loopback =-466;
27120: waveform_sig_loopback =-312;
27121: waveform_sig_loopback =-2318;
27122: waveform_sig_loopback =-82;
27123: waveform_sig_loopback =-836;
27124: waveform_sig_loopback =-1750;
27125: waveform_sig_loopback =-1120;
27126: waveform_sig_loopback =-439;
27127: waveform_sig_loopback =-1539;
27128: waveform_sig_loopback =-2169;
27129: waveform_sig_loopback =-278;
27130: waveform_sig_loopback =-913;
27131: waveform_sig_loopback =-3178;
27132: waveform_sig_loopback =-684;
27133: waveform_sig_loopback =-179;
27134: waveform_sig_loopback =-3102;
27135: waveform_sig_loopback =-1861;
27136: waveform_sig_loopback =-62;
27137: waveform_sig_loopback =-2670;
27138: waveform_sig_loopback =-874;
27139: waveform_sig_loopback =-1492;
27140: waveform_sig_loopback =-5026;
27141: waveform_sig_loopback =437;
27142: waveform_sig_loopback =-1015;
27143: waveform_sig_loopback =-2605;
27144: waveform_sig_loopback =-3130;
27145: waveform_sig_loopback =-2350;
27146: waveform_sig_loopback =-206;
27147: waveform_sig_loopback =-2099;
27148: waveform_sig_loopback =-3789;
27149: waveform_sig_loopback =-1241;
27150: waveform_sig_loopback =-2640;
27151: waveform_sig_loopback =-1798;
27152: waveform_sig_loopback =-2555;
27153: waveform_sig_loopback =-3327;
27154: waveform_sig_loopback =-773;
27155: waveform_sig_loopback =-3464;
27156: waveform_sig_loopback =-2542;
27157: waveform_sig_loopback =-2211;
27158: waveform_sig_loopback =-2711;
27159: waveform_sig_loopback =-3131;
27160: waveform_sig_loopback =-2105;
27161: waveform_sig_loopback =-2501;
27162: waveform_sig_loopback =-3839;
27163: waveform_sig_loopback =-1990;
27164: waveform_sig_loopback =-2818;
27165: waveform_sig_loopback =-3200;
27166: waveform_sig_loopback =-3438;
27167: waveform_sig_loopback =-1772;
27168: waveform_sig_loopback =-3536;
27169: waveform_sig_loopback =-4187;
27170: waveform_sig_loopback =-1461;
27171: waveform_sig_loopback =-3373;
27172: waveform_sig_loopback =-4630;
27173: waveform_sig_loopback =-2303;
27174: waveform_sig_loopback =-2436;
27175: waveform_sig_loopback =-4447;
27176: waveform_sig_loopback =-3912;
27177: waveform_sig_loopback =-1791;
27178: waveform_sig_loopback =-4358;
27179: waveform_sig_loopback =-2778;
27180: waveform_sig_loopback =-3261;
27181: waveform_sig_loopback =-6775;
27182: waveform_sig_loopback =-1188;
27183: waveform_sig_loopback =-2781;
27184: waveform_sig_loopback =-4482;
27185: waveform_sig_loopback =-4835;
27186: waveform_sig_loopback =-3860;
27187: waveform_sig_loopback =-2004;
27188: waveform_sig_loopback =-4017;
27189: waveform_sig_loopback =-5248;
27190: waveform_sig_loopback =-3035;
27191: waveform_sig_loopback =-4399;
27192: waveform_sig_loopback =-3326;
27193: waveform_sig_loopback =-4534;
27194: waveform_sig_loopback =-4671;
27195: waveform_sig_loopback =-2593;
27196: waveform_sig_loopback =-5352;
27197: waveform_sig_loopback =-3857;
27198: waveform_sig_loopback =-4077;
27199: waveform_sig_loopback =-4342;
27200: waveform_sig_loopback =-4622;
27201: waveform_sig_loopback =-4039;
27202: waveform_sig_loopback =-3901;
27203: waveform_sig_loopback =-5499;
27204: waveform_sig_loopback =-3900;
27205: waveform_sig_loopback =-4060;
27206: waveform_sig_loopback =-5224;
27207: waveform_sig_loopback =-4844;
27208: waveform_sig_loopback =-3294;
27209: waveform_sig_loopback =-5606;
27210: waveform_sig_loopback =-5348;
27211: waveform_sig_loopback =-3199;
27212: waveform_sig_loopback =-5163;
27213: waveform_sig_loopback =-5950;
27214: waveform_sig_loopback =-3996;
27215: waveform_sig_loopback =-3982;
27216: waveform_sig_loopback =-5971;
27217: waveform_sig_loopback =-5555;
27218: waveform_sig_loopback =-3134;
27219: waveform_sig_loopback =-6020;
27220: waveform_sig_loopback =-4256;
27221: waveform_sig_loopback =-4809;
27222: waveform_sig_loopback =-8272;
27223: waveform_sig_loopback =-2608;
27224: waveform_sig_loopback =-4316;
27225: waveform_sig_loopback =-6131;
27226: waveform_sig_loopback =-6252;
27227: waveform_sig_loopback =-5090;
27228: waveform_sig_loopback =-3712;
27229: waveform_sig_loopback =-5483;
27230: waveform_sig_loopback =-6545;
27231: waveform_sig_loopback =-4658;
27232: waveform_sig_loopback =-5572;
27233: waveform_sig_loopback =-4932;
27234: waveform_sig_loopback =-6029;
27235: waveform_sig_loopback =-5690;
27236: waveform_sig_loopback =-4386;
27237: waveform_sig_loopback =-6503;
27238: waveform_sig_loopback =-5170;
27239: waveform_sig_loopback =-5772;
27240: waveform_sig_loopback =-5257;
27241: waveform_sig_loopback =-6319;
27242: waveform_sig_loopback =-5216;
27243: waveform_sig_loopback =-5153;
27244: waveform_sig_loopback =-7217;
27245: waveform_sig_loopback =-4760;
27246: waveform_sig_loopback =-5510;
27247: waveform_sig_loopback =-6680;
27248: waveform_sig_loopback =-5736;
27249: waveform_sig_loopback =-4911;
27250: waveform_sig_loopback =-6719;
27251: waveform_sig_loopback =-6467;
27252: waveform_sig_loopback =-4541;
27253: waveform_sig_loopback =-6404;
27254: waveform_sig_loopback =-7163;
27255: waveform_sig_loopback =-5146;
27256: waveform_sig_loopback =-5243;
27257: waveform_sig_loopback =-7214;
27258: waveform_sig_loopback =-6764;
27259: waveform_sig_loopback =-4142;
27260: waveform_sig_loopback =-7408;
27261: waveform_sig_loopback =-5303;
27262: waveform_sig_loopback =-5978;
27263: waveform_sig_loopback =-9603;
27264: waveform_sig_loopback =-3447;
27265: waveform_sig_loopback =-5544;
27266: waveform_sig_loopback =-7462;
27267: waveform_sig_loopback =-7081;
27268: waveform_sig_loopback =-6354;
27269: waveform_sig_loopback =-4782;
27270: waveform_sig_loopback =-6365;
27271: waveform_sig_loopback =-7990;
27272: waveform_sig_loopback =-5425;
27273: waveform_sig_loopback =-6637;
27274: waveform_sig_loopback =-6184;
27275: waveform_sig_loopback =-6773;
27276: waveform_sig_loopback =-6949;
27277: waveform_sig_loopback =-5347;
27278: waveform_sig_loopback =-7368;
27279: waveform_sig_loopback =-6407;
27280: waveform_sig_loopback =-6574;
27281: waveform_sig_loopback =-6283;
27282: waveform_sig_loopback =-7404;
27283: waveform_sig_loopback =-5888;
27284: waveform_sig_loopback =-6333;
27285: waveform_sig_loopback =-8105;
27286: waveform_sig_loopback =-5435;
27287: waveform_sig_loopback =-6733;
27288: waveform_sig_loopback =-7489;
27289: waveform_sig_loopback =-6438;
27290: waveform_sig_loopback =-6003;
27291: waveform_sig_loopback =-7532;
27292: waveform_sig_loopback =-7252;
27293: waveform_sig_loopback =-5534;
27294: waveform_sig_loopback =-7079;
27295: waveform_sig_loopback =-8114;
27296: waveform_sig_loopback =-5934;
27297: waveform_sig_loopback =-5911;
27298: waveform_sig_loopback =-8389;
27299: waveform_sig_loopback =-7424;
27300: waveform_sig_loopback =-4762;
27301: waveform_sig_loopback =-8457;
27302: waveform_sig_loopback =-5643;
27303: waveform_sig_loopback =-7364;
27304: waveform_sig_loopback =-10056;
27305: waveform_sig_loopback =-3642;
27306: waveform_sig_loopback =-6857;
27307: waveform_sig_loopback =-8071;
27308: waveform_sig_loopback =-7677;
27309: waveform_sig_loopback =-7073;
27310: waveform_sig_loopback =-5240;
27311: waveform_sig_loopback =-7465;
27312: waveform_sig_loopback =-8535;
27313: waveform_sig_loopback =-5772;
27314: waveform_sig_loopback =-7632;
27315: waveform_sig_loopback =-6700;
27316: waveform_sig_loopback =-7370;
27317: waveform_sig_loopback =-7555;
27318: waveform_sig_loopback =-5873;
27319: waveform_sig_loopback =-8090;
27320: waveform_sig_loopback =-7033;
27321: waveform_sig_loopback =-6812;
27322: waveform_sig_loopback =-7153;
27323: waveform_sig_loopback =-7982;
27324: waveform_sig_loopback =-6095;
27325: waveform_sig_loopback =-7248;
27326: waveform_sig_loopback =-8300;
27327: waveform_sig_loopback =-6025;
27328: waveform_sig_loopback =-7390;
27329: waveform_sig_loopback =-7633;
27330: waveform_sig_loopback =-7175;
27331: waveform_sig_loopback =-6413;
27332: waveform_sig_loopback =-7881;
27333: waveform_sig_loopback =-7808;
27334: waveform_sig_loopback =-5818;
27335: waveform_sig_loopback =-7565;
27336: waveform_sig_loopback =-8530;
27337: waveform_sig_loopback =-6064;
27338: waveform_sig_loopback =-6421;
27339: waveform_sig_loopback =-8770;
27340: waveform_sig_loopback =-7213;
27341: waveform_sig_loopback =-5460;
27342: waveform_sig_loopback =-8856;
27343: waveform_sig_loopback =-5522;
27344: waveform_sig_loopback =-8037;
27345: waveform_sig_loopback =-10001;
27346: waveform_sig_loopback =-4034;
27347: waveform_sig_loopback =-7354;
27348: waveform_sig_loopback =-7787;
27349: waveform_sig_loopback =-8325;
27350: waveform_sig_loopback =-7224;
27351: waveform_sig_loopback =-5157;
27352: waveform_sig_loopback =-8085;
27353: waveform_sig_loopback =-8298;
27354: waveform_sig_loopback =-6119;
27355: waveform_sig_loopback =-7932;
27356: waveform_sig_loopback =-6373;
27357: waveform_sig_loopback =-7951;
27358: waveform_sig_loopback =-7510;
27359: waveform_sig_loopback =-5814;
27360: waveform_sig_loopback =-8423;
27361: waveform_sig_loopback =-6868;
27362: waveform_sig_loopback =-7022;
27363: waveform_sig_loopback =-7269;
27364: waveform_sig_loopback =-7735;
27365: waveform_sig_loopback =-6292;
27366: waveform_sig_loopback =-7432;
27367: waveform_sig_loopback =-7927;
27368: waveform_sig_loopback =-6255;
27369: waveform_sig_loopback =-7309;
27370: waveform_sig_loopback =-7551;
27371: waveform_sig_loopback =-7269;
27372: waveform_sig_loopback =-6074;
27373: waveform_sig_loopback =-8074;
27374: waveform_sig_loopback =-7670;
27375: waveform_sig_loopback =-5513;
27376: waveform_sig_loopback =-7798;
27377: waveform_sig_loopback =-8285;
27378: waveform_sig_loopback =-5818;
27379: waveform_sig_loopback =-6534;
27380: waveform_sig_loopback =-8536;
27381: waveform_sig_loopback =-6927;
27382: waveform_sig_loopback =-5548;
27383: waveform_sig_loopback =-8436;
27384: waveform_sig_loopback =-5298;
27385: waveform_sig_loopback =-8223;
27386: waveform_sig_loopback =-9263;
27387: waveform_sig_loopback =-4069;
27388: waveform_sig_loopback =-7072;
27389: waveform_sig_loopback =-7421;
27390: waveform_sig_loopback =-8362;
27391: waveform_sig_loopback =-6421;
27392: waveform_sig_loopback =-5115;
27393: waveform_sig_loopback =-7953;
27394: waveform_sig_loopback =-7565;
27395: waveform_sig_loopback =-6187;
27396: waveform_sig_loopback =-7303;
27397: waveform_sig_loopback =-6041;
27398: waveform_sig_loopback =-7904;
27399: waveform_sig_loopback =-6615;
27400: waveform_sig_loopback =-5810;
27401: waveform_sig_loopback =-7956;
27402: waveform_sig_loopback =-6269;
27403: waveform_sig_loopback =-6799;
27404: waveform_sig_loopback =-6679;
27405: waveform_sig_loopback =-7373;
27406: waveform_sig_loopback =-5790;
27407: waveform_sig_loopback =-6957;
27408: waveform_sig_loopback =-7404;
27409: waveform_sig_loopback =-5825;
27410: waveform_sig_loopback =-6708;
27411: waveform_sig_loopback =-7053;
27412: waveform_sig_loopback =-6756;
27413: waveform_sig_loopback =-5357;
27414: waveform_sig_loopback =-7793;
27415: waveform_sig_loopback =-6904;
27416: waveform_sig_loopback =-4780;
27417: waveform_sig_loopback =-7618;
27418: waveform_sig_loopback =-7317;
27419: waveform_sig_loopback =-5243;
27420: waveform_sig_loopback =-6167;
27421: waveform_sig_loopback =-7572;
27422: waveform_sig_loopback =-6557;
27423: waveform_sig_loopback =-4784;
27424: waveform_sig_loopback =-7659;
27425: waveform_sig_loopback =-4910;
27426: waveform_sig_loopback =-7298;
27427: waveform_sig_loopback =-8571;
27428: waveform_sig_loopback =-3380;
27429: waveform_sig_loopback =-6094;
27430: waveform_sig_loopback =-7185;
27431: waveform_sig_loopback =-7250;
27432: waveform_sig_loopback =-5631;
27433: waveform_sig_loopback =-4666;
27434: waveform_sig_loopback =-6838;
27435: waveform_sig_loopback =-7007;
27436: waveform_sig_loopback =-5327;
27437: waveform_sig_loopback =-6385;
27438: waveform_sig_loopback =-5427;
27439: waveform_sig_loopback =-6910;
27440: waveform_sig_loopback =-5739;
27441: waveform_sig_loopback =-5115;
27442: waveform_sig_loopback =-6974;
27443: waveform_sig_loopback =-5384;
27444: waveform_sig_loopback =-6005;
27445: waveform_sig_loopback =-5746;
27446: waveform_sig_loopback =-6402;
27447: waveform_sig_loopback =-4987;
27448: waveform_sig_loopback =-5864;
27449: waveform_sig_loopback =-6586;
27450: waveform_sig_loopback =-4883;
27451: waveform_sig_loopback =-5474;
27452: waveform_sig_loopback =-6574;
27453: waveform_sig_loopback =-5285;
27454: waveform_sig_loopback =-4576;
27455: waveform_sig_loopback =-7015;
27456: waveform_sig_loopback =-5325;
27457: waveform_sig_loopback =-4315;
27458: waveform_sig_loopback =-6352;
27459: waveform_sig_loopback =-6134;
27460: waveform_sig_loopback =-4478;
27461: waveform_sig_loopback =-4778;
27462: waveform_sig_loopback =-6805;
27463: waveform_sig_loopback =-5310;
27464: waveform_sig_loopback =-3534;
27465: waveform_sig_loopback =-6934;
27466: waveform_sig_loopback =-3474;
27467: waveform_sig_loopback =-6402;
27468: waveform_sig_loopback =-7466;
27469: waveform_sig_loopback =-1980;
27470: waveform_sig_loopback =-5215;
27471: waveform_sig_loopback =-6092;
27472: waveform_sig_loopback =-5825;
27473: waveform_sig_loopback =-4604;
27474: waveform_sig_loopback =-3412;
27475: waveform_sig_loopback =-5649;
27476: waveform_sig_loopback =-5885;
27477: waveform_sig_loopback =-3900;
27478: waveform_sig_loopback =-5193;
27479: waveform_sig_loopback =-4270;
27480: waveform_sig_loopback =-5550;
27481: waveform_sig_loopback =-4449;
27482: waveform_sig_loopback =-3963;
27483: waveform_sig_loopback =-5556;
27484: waveform_sig_loopback =-4166;
27485: waveform_sig_loopback =-4731;
27486: waveform_sig_loopback =-4229;
27487: waveform_sig_loopback =-5351;
27488: waveform_sig_loopback =-3453;
27489: waveform_sig_loopback =-4562;
27490: waveform_sig_loopback =-5491;
27491: waveform_sig_loopback =-3079;
27492: waveform_sig_loopback =-4551;
27493: waveform_sig_loopback =-5115;
27494: waveform_sig_loopback =-3506;
27495: waveform_sig_loopback =-3788;
27496: waveform_sig_loopback =-5179;
27497: waveform_sig_loopback =-4020;
27498: waveform_sig_loopback =-3056;
27499: waveform_sig_loopback =-4612;
27500: waveform_sig_loopback =-5091;
27501: waveform_sig_loopback =-2658;
27502: waveform_sig_loopback =-3461;
27503: waveform_sig_loopback =-5572;
27504: waveform_sig_loopback =-3363;
27505: waveform_sig_loopback =-2389;
27506: waveform_sig_loopback =-5359;
27507: waveform_sig_loopback =-1796;
27508: waveform_sig_loopback =-5323;
27509: waveform_sig_loopback =-5567;
27510: waveform_sig_loopback =-504;
27511: waveform_sig_loopback =-3817;
27512: waveform_sig_loopback =-4496;
27513: waveform_sig_loopback =-4266;
27514: waveform_sig_loopback =-3082;
27515: waveform_sig_loopback =-1761;
27516: waveform_sig_loopback =-4193;
27517: waveform_sig_loopback =-4424;
27518: waveform_sig_loopback =-2126;
27519: waveform_sig_loopback =-3789;
27520: waveform_sig_loopback =-2663;
27521: waveform_sig_loopback =-3874;
27522: waveform_sig_loopback =-3055;
27523: waveform_sig_loopback =-2201;
27524: waveform_sig_loopback =-3971;
27525: waveform_sig_loopback =-2769;
27526: waveform_sig_loopback =-2759;
27527: waveform_sig_loopback =-2957;
27528: waveform_sig_loopback =-3631;
27529: waveform_sig_loopback =-1521;
27530: waveform_sig_loopback =-3513;
27531: waveform_sig_loopback =-3317;
27532: waveform_sig_loopback =-1626;
27533: waveform_sig_loopback =-3053;
27534: waveform_sig_loopback =-3142;
27535: waveform_sig_loopback =-2182;
27536: waveform_sig_loopback =-1886;
27537: waveform_sig_loopback =-3566;
27538: waveform_sig_loopback =-2358;
27539: waveform_sig_loopback =-1240;
27540: waveform_sig_loopback =-3087;
27541: waveform_sig_loopback =-3334;
27542: waveform_sig_loopback =-897;
27543: waveform_sig_loopback =-1809;
27544: waveform_sig_loopback =-4003;
27545: waveform_sig_loopback =-1341;
27546: waveform_sig_loopback =-935;
27547: waveform_sig_loopback =-3614;
27548: waveform_sig_loopback =220;
27549: waveform_sig_loopback =-4190;
27550: waveform_sig_loopback =-3315;
27551: waveform_sig_loopback =1220;
27552: waveform_sig_loopback =-2393;
27553: waveform_sig_loopback =-2389;
27554: waveform_sig_loopback =-2750;
27555: waveform_sig_loopback =-1166;
27556: waveform_sig_loopback =198;
27557: waveform_sig_loopback =-2897;
27558: waveform_sig_loopback =-2257;
27559: waveform_sig_loopback =-418;
27560: waveform_sig_loopback =-2209;
27561: waveform_sig_loopback =-476;
27562: waveform_sig_loopback =-2467;
27563: waveform_sig_loopback =-1031;
27564: waveform_sig_loopback =-292;
27565: waveform_sig_loopback =-2471;
27566: waveform_sig_loopback =-659;
27567: waveform_sig_loopback =-1074;
27568: waveform_sig_loopback =-1267;
27569: waveform_sig_loopback =-1555;
27570: waveform_sig_loopback =99;
27571: waveform_sig_loopback =-1731;
27572: waveform_sig_loopback =-1284;
27573: waveform_sig_loopback =39;
27574: waveform_sig_loopback =-1134;
27575: waveform_sig_loopback =-1265;
27576: waveform_sig_loopback =-399;
27577: waveform_sig_loopback =25;
27578: waveform_sig_loopback =-1749;
27579: waveform_sig_loopback =-597;
27580: waveform_sig_loopback =797;
27581: waveform_sig_loopback =-1457;
27582: waveform_sig_loopback =-1386;
27583: waveform_sig_loopback =1229;
27584: waveform_sig_loopback =-345;
27585: waveform_sig_loopback =-1897;
27586: waveform_sig_loopback =662;
27587: waveform_sig_loopback =574;
27588: waveform_sig_loopback =-1373;
27589: waveform_sig_loopback =1941;
27590: waveform_sig_loopback =-2505;
27591: waveform_sig_loopback =-865;
27592: waveform_sig_loopback =2623;
27593: waveform_sig_loopback =-358;
27594: waveform_sig_loopback =-435;
27595: waveform_sig_loopback =-1147;
27596: waveform_sig_loopback =1165;
27597: waveform_sig_loopback =1812;
27598: waveform_sig_loopback =-1078;
27599: waveform_sig_loopback =37;
27600: waveform_sig_loopback =1005;
27601: waveform_sig_loopback =57;
27602: waveform_sig_loopback =1387;
27603: waveform_sig_loopback =-886;
27604: waveform_sig_loopback =1327;
27605: waveform_sig_loopback =1310;
27606: waveform_sig_loopback =-517;
27607: waveform_sig_loopback =1419;
27608: waveform_sig_loopback =611;
27609: waveform_sig_loopback =787;
27610: waveform_sig_loopback =403;
27611: waveform_sig_loopback =1907;
27612: waveform_sig_loopback =186;
27613: waveform_sig_loopback =777;
27614: waveform_sig_loopback =1765;
27615: waveform_sig_loopback =952;
27616: waveform_sig_loopback =512;
27617: waveform_sig_loopback =1530;
27618: waveform_sig_loopback =2163;
27619: waveform_sig_loopback =-255;
27620: waveform_sig_loopback =1656;
27621: waveform_sig_loopback =2745;
27622: waveform_sig_loopback =66;
27623: waveform_sig_loopback =967;
27624: waveform_sig_loopback =2915;
27625: waveform_sig_loopback =1445;
27626: waveform_sig_loopback =291;
27627: waveform_sig_loopback =2244;
27628: waveform_sig_loopback =2675;
27629: waveform_sig_loopback =558;
27630: waveform_sig_loopback =3587;
27631: waveform_sig_loopback =-439;
27632: waveform_sig_loopback =912;
27633: waveform_sig_loopback =4637;
27634: waveform_sig_loopback =1634;
27635: waveform_sig_loopback =1042;
27636: waveform_sig_loopback =1071;
27637: waveform_sig_loopback =3088;
27638: waveform_sig_loopback =3467;
27639: waveform_sig_loopback =922;
27640: waveform_sig_loopback =1878;
27641: waveform_sig_loopback =2889;
27642: waveform_sig_loopback =1925;
27643: waveform_sig_loopback =3054;
27644: waveform_sig_loopback =1060;
27645: waveform_sig_loopback =3317;
27646: waveform_sig_loopback =2812;
27647: waveform_sig_loopback =1273;
27648: waveform_sig_loopback =3455;
27649: waveform_sig_loopback =2285;
27650: waveform_sig_loopback =2751;
27651: waveform_sig_loopback =2041;
27652: waveform_sig_loopback =3605;
27653: waveform_sig_loopback =2504;
27654: waveform_sig_loopback =2142;
27655: waveform_sig_loopback =3693;
27656: waveform_sig_loopback =2757;
27657: waveform_sig_loopback =2195;
27658: waveform_sig_loopback =3786;
27659: waveform_sig_loopback =3377;
27660: waveform_sig_loopback =1712;
27661: waveform_sig_loopback =3757;
27662: waveform_sig_loopback =4129;
27663: waveform_sig_loopback =1916;
27664: waveform_sig_loopback =2834;
27665: waveform_sig_loopback =4661;
27666: waveform_sig_loopback =3196;
27667: waveform_sig_loopback =1929;
27668: waveform_sig_loopback =4127;
27669: waveform_sig_loopback =4506;
27670: waveform_sig_loopback =2144;
27671: waveform_sig_loopback =5413;
27672: waveform_sig_loopback =1249;
27673: waveform_sig_loopback =2698;
27674: waveform_sig_loopback =6446;
27675: waveform_sig_loopback =3193;
27676: waveform_sig_loopback =2658;
27677: waveform_sig_loopback =3086;
27678: waveform_sig_loopback =4628;
27679: waveform_sig_loopback =5065;
27680: waveform_sig_loopback =2761;
27681: waveform_sig_loopback =3464;
27682: waveform_sig_loopback =4643;
27683: waveform_sig_loopback =3711;
27684: waveform_sig_loopback =4548;
27685: waveform_sig_loopback =3010;
27686: waveform_sig_loopback =4921;
27687: waveform_sig_loopback =4313;
27688: waveform_sig_loopback =3488;
27689: waveform_sig_loopback =4637;
27690: waveform_sig_loopback =4042;
27691: waveform_sig_loopback =4511;
27692: waveform_sig_loopback =3539;
27693: waveform_sig_loopback =5632;
27694: waveform_sig_loopback =3613;
27695: waveform_sig_loopback =3870;
27696: waveform_sig_loopback =5665;
27697: waveform_sig_loopback =3980;
27698: waveform_sig_loopback =3836;
27699: waveform_sig_loopback =5435;
27700: waveform_sig_loopback =4814;
27701: waveform_sig_loopback =3467;
27702: waveform_sig_loopback =5177;
27703: waveform_sig_loopback =5610;
27704: waveform_sig_loopback =3673;
27705: waveform_sig_loopback =4283;
27706: waveform_sig_loopback =6176;
27707: waveform_sig_loopback =4823;
27708: waveform_sig_loopback =3369;
27709: waveform_sig_loopback =5837;
27710: waveform_sig_loopback =5885;
27711: waveform_sig_loopback =3586;
27712: waveform_sig_loopback =7164;
27713: waveform_sig_loopback =2362;
27714: waveform_sig_loopback =4325;
27715: waveform_sig_loopback =8185;
27716: waveform_sig_loopback =4291;
27717: waveform_sig_loopback =4190;
27718: waveform_sig_loopback =4632;
27719: waveform_sig_loopback =5904;
27720: waveform_sig_loopback =6794;
27721: waveform_sig_loopback =3916;
27722: waveform_sig_loopback =4863;
27723: waveform_sig_loopback =6263;
27724: waveform_sig_loopback =4867;
27725: waveform_sig_loopback =5986;
27726: waveform_sig_loopback =4470;
27727: waveform_sig_loopback =6172;
27728: waveform_sig_loopback =5836;
27729: waveform_sig_loopback =4821;
27730: waveform_sig_loopback =5890;
27731: waveform_sig_loopback =5702;
27732: waveform_sig_loopback =5499;
27733: waveform_sig_loopback =5079;
27734: waveform_sig_loopback =7081;
27735: waveform_sig_loopback =4558;
27736: waveform_sig_loopback =5607;
27737: waveform_sig_loopback =6780;
27738: waveform_sig_loopback =5202;
27739: waveform_sig_loopback =5361;
27740: waveform_sig_loopback =6635;
27741: waveform_sig_loopback =6044;
27742: waveform_sig_loopback =4818;
27743: waveform_sig_loopback =6477;
27744: waveform_sig_loopback =6809;
27745: waveform_sig_loopback =4949;
27746: waveform_sig_loopback =5410;
27747: waveform_sig_loopback =7550;
27748: waveform_sig_loopback =5923;
27749: waveform_sig_loopback =4364;
27750: waveform_sig_loopback =7496;
27751: waveform_sig_loopback =6626;
27752: waveform_sig_loopback =4917;
27753: waveform_sig_loopback =8533;
27754: waveform_sig_loopback =2918;
27755: waveform_sig_loopback =6207;
27756: waveform_sig_loopback =8986;
27757: waveform_sig_loopback =5203;
27758: waveform_sig_loopback =5734;
27759: waveform_sig_loopback =5364;
27760: waveform_sig_loopback =7289;
27761: waveform_sig_loopback =7856;
27762: waveform_sig_loopback =4633;
27763: waveform_sig_loopback =6401;
27764: waveform_sig_loopback =7114;
27765: waveform_sig_loopback =5939;
27766: waveform_sig_loopback =7186;
27767: waveform_sig_loopback =5256;
27768: waveform_sig_loopback =7368;
27769: waveform_sig_loopback =6836;
27770: waveform_sig_loopback =5642;
27771: waveform_sig_loopback =6995;
27772: waveform_sig_loopback =6742;
27773: waveform_sig_loopback =6255;
27774: waveform_sig_loopback =6288;
27775: waveform_sig_loopback =7934;
27776: waveform_sig_loopback =5335;
27777: waveform_sig_loopback =6899;
27778: waveform_sig_loopback =7390;
27779: waveform_sig_loopback =6170;
27780: waveform_sig_loopback =6445;
27781: waveform_sig_loopback =7245;
27782: waveform_sig_loopback =7185;
27783: waveform_sig_loopback =5540;
27784: waveform_sig_loopback =7353;
27785: waveform_sig_loopback =7894;
27786: waveform_sig_loopback =5393;
27787: waveform_sig_loopback =6582;
27788: waveform_sig_loopback =8441;
27789: waveform_sig_loopback =6425;
27790: waveform_sig_loopback =5406;
27791: waveform_sig_loopback =8324;
27792: waveform_sig_loopback =7162;
27793: waveform_sig_loopback =5973;
27794: waveform_sig_loopback =9126;
27795: waveform_sig_loopback =3482;
27796: waveform_sig_loopback =7474;
27797: waveform_sig_loopback =9345;
27798: waveform_sig_loopback =5995;
27799: waveform_sig_loopback =6536;
27800: waveform_sig_loopback =5837;
27801: waveform_sig_loopback =8380;
27802: waveform_sig_loopback =8248;
27803: waveform_sig_loopback =5162;
27804: waveform_sig_loopback =7495;
27805: waveform_sig_loopback =7311;
27806: waveform_sig_loopback =6802;
27807: waveform_sig_loopback =7806;
27808: waveform_sig_loopback =5617;
27809: waveform_sig_loopback =8374;
27810: waveform_sig_loopback =7089;
27811: waveform_sig_loopback =6269;
27812: waveform_sig_loopback =7780;
27813: waveform_sig_loopback =7015;
27814: waveform_sig_loopback =6906;
27815: waveform_sig_loopback =6922;
27816: waveform_sig_loopback =8194;
27817: waveform_sig_loopback =5995;
27818: waveform_sig_loopback =7407;
27819: waveform_sig_loopback =7743;
27820: waveform_sig_loopback =6804;
27821: waveform_sig_loopback =6737;
27822: waveform_sig_loopback =7789;
27823: waveform_sig_loopback =7651;
27824: waveform_sig_loopback =5766;
27825: waveform_sig_loopback =7968;
27826: waveform_sig_loopback =8244;
27827: waveform_sig_loopback =5583;
27828: waveform_sig_loopback =7189;
27829: waveform_sig_loopback =8667;
27830: waveform_sig_loopback =6556;
27831: waveform_sig_loopback =6138;
27832: waveform_sig_loopback =8360;
27833: waveform_sig_loopback =7486;
27834: waveform_sig_loopback =6543;
27835: waveform_sig_loopback =9013;
27836: waveform_sig_loopback =3968;
27837: waveform_sig_loopback =7774;
27838: waveform_sig_loopback =9494;
27839: waveform_sig_loopback =6414;
27840: waveform_sig_loopback =6464;
27841: waveform_sig_loopback =6253;
27842: waveform_sig_loopback =8767;
27843: waveform_sig_loopback =8098;
27844: waveform_sig_loopback =5529;
27845: waveform_sig_loopback =7700;
27846: waveform_sig_loopback =7201;
27847: waveform_sig_loopback =7367;
27848: waveform_sig_loopback =7512;
27849: waveform_sig_loopback =5892;
27850: waveform_sig_loopback =8696;
27851: waveform_sig_loopback =6691;
27852: waveform_sig_loopback =6810;
27853: waveform_sig_loopback =7612;
27854: waveform_sig_loopback =7062;
27855: waveform_sig_loopback =7106;
27856: waveform_sig_loopback =6777;
27857: waveform_sig_loopback =8364;
27858: waveform_sig_loopback =5919;
27859: waveform_sig_loopback =7395;
27860: waveform_sig_loopback =7770;
27861: waveform_sig_loopback =6766;
27862: waveform_sig_loopback =6619;
27863: waveform_sig_loopback =7878;
27864: waveform_sig_loopback =7464;
27865: waveform_sig_loopback =5569;
27866: waveform_sig_loopback =8199;
27867: waveform_sig_loopback =7855;
27868: waveform_sig_loopback =5407;
27869: waveform_sig_loopback =7461;
27870: waveform_sig_loopback =8208;
27871: waveform_sig_loopback =6563;
27872: waveform_sig_loopback =5936;
27873: waveform_sig_loopback =8135;
27874: waveform_sig_loopback =7512;
27875: waveform_sig_loopback =6128;
27876: waveform_sig_loopback =8808;
27877: waveform_sig_loopback =3870;
27878: waveform_sig_loopback =7399;
27879: waveform_sig_loopback =9398;
27880: waveform_sig_loopback =6057;
27881: waveform_sig_loopback =5960;
27882: waveform_sig_loopback =6471;
27883: waveform_sig_loopback =8053;
27884: waveform_sig_loopback =7872;
27885: waveform_sig_loopback =5365;
27886: waveform_sig_loopback =7112;
27887: waveform_sig_loopback =7165;
27888: waveform_sig_loopback =6811;
27889: waveform_sig_loopback =7124;
27890: waveform_sig_loopback =5799;
27891: waveform_sig_loopback =8037;
27892: waveform_sig_loopback =6417;
27893: waveform_sig_loopback =6385;
27894: waveform_sig_loopback =7181;
27895: waveform_sig_loopback =6672;
27896: waveform_sig_loopback =6580;
27897: waveform_sig_loopback =6502;
27898: waveform_sig_loopback =7747;
27899: waveform_sig_loopback =5626;
27900: waveform_sig_loopback =6698;
27901: waveform_sig_loopback =7446;
27902: waveform_sig_loopback =6245;
27903: waveform_sig_loopback =5853;
27904: waveform_sig_loopback =7864;
27905: waveform_sig_loopback =6340;
27906: waveform_sig_loopback =5357;
27907: waveform_sig_loopback =7756;
27908: waveform_sig_loopback =6751;
27909: waveform_sig_loopback =5389;
27910: waveform_sig_loopback =6486;
27911: waveform_sig_loopback =7629;
27912: waveform_sig_loopback =6156;
27913: waveform_sig_loopback =4870;
27914: waveform_sig_loopback =8051;
27915: waveform_sig_loopback =6408;
27916: waveform_sig_loopback =5513;
27917: waveform_sig_loopback =8413;
27918: waveform_sig_loopback =2658;
27919: waveform_sig_loopback =7262;
27920: waveform_sig_loopback =8512;
27921: waveform_sig_loopback =5065;
27922: waveform_sig_loopback =5503;
27923: waveform_sig_loopback =5600;
27924: waveform_sig_loopback =7359;
27925: waveform_sig_loopback =7092;
27926: waveform_sig_loopback =4488;
27927: waveform_sig_loopback =6397;
27928: waveform_sig_loopback =6397;
27929: waveform_sig_loopback =5893;
27930: waveform_sig_loopback =6302;
27931: waveform_sig_loopback =5039;
27932: waveform_sig_loopback =7052;
27933: waveform_sig_loopback =5596;
27934: waveform_sig_loopback =5590;
27935: waveform_sig_loopback =6119;
27936: waveform_sig_loopback =5938;
27937: waveform_sig_loopback =5595;
27938: waveform_sig_loopback =5445;
27939: waveform_sig_loopback =7141;
27940: waveform_sig_loopback =4311;
27941: waveform_sig_loopback =5977;
27942: waveform_sig_loopback =6598;
27943: waveform_sig_loopback =4778;
27944: waveform_sig_loopback =5537;
27945: waveform_sig_loopback =6489;
27946: waveform_sig_loopback =5230;
27947: waveform_sig_loopback =4740;
27948: waveform_sig_loopback =6355;
27949: waveform_sig_loopback =6011;
27950: waveform_sig_loopback =4262;
27951: waveform_sig_loopback =5296;
27952: waveform_sig_loopback =7032;
27953: waveform_sig_loopback =4602;
27954: waveform_sig_loopback =3961;
27955: waveform_sig_loopback =7231;
27956: waveform_sig_loopback =4808;
27957: waveform_sig_loopback =4953;
27958: waveform_sig_loopback =6924;
27959: waveform_sig_loopback =1481;
27960: waveform_sig_loopback =6584;
27961: waveform_sig_loopback =6949;
27962: waveform_sig_loopback =4150;
27963: waveform_sig_loopback =4237;
27964: waveform_sig_loopback =4446;
27965: waveform_sig_loopback =6277;
27966: waveform_sig_loopback =5818;
27967: waveform_sig_loopback =3228;
27968: waveform_sig_loopback =5180;
27969: waveform_sig_loopback =5275;
27970: waveform_sig_loopback =4548;
27971: waveform_sig_loopback =5140;
27972: waveform_sig_loopback =3761;
27973: waveform_sig_loopback =5752;
27974: waveform_sig_loopback =4574;
27975: waveform_sig_loopback =4092;
27976: waveform_sig_loopback =4857;
27977: waveform_sig_loopback =4917;
27978: waveform_sig_loopback =3822;
27979: waveform_sig_loopback =4693;
27980: waveform_sig_loopback =5500;
27981: waveform_sig_loopback =2783;
27982: waveform_sig_loopback =5280;
27983: waveform_sig_loopback =4606;
27984: waveform_sig_loopback =3837;
27985: waveform_sig_loopback =4049;
27986: waveform_sig_loopback =4951;
27987: waveform_sig_loopback =4281;
27988: waveform_sig_loopback =2934;
27989: waveform_sig_loopback =5214;
27990: waveform_sig_loopback =4618;
27991: waveform_sig_loopback =2505;
27992: waveform_sig_loopback =4302;
27993: waveform_sig_loopback =5365;
27994: waveform_sig_loopback =3108;
27995: waveform_sig_loopback =2540;
27996: waveform_sig_loopback =5684;
27997: waveform_sig_loopback =3413;
27998: waveform_sig_loopback =3603;
27999: waveform_sig_loopback =5209;
28000: waveform_sig_loopback =-255;
28001: waveform_sig_loopback =5659;
28002: waveform_sig_loopback =5244;
28003: waveform_sig_loopback =2383;
28004: waveform_sig_loopback =2889;
28005: waveform_sig_loopback =2832;
28006: waveform_sig_loopback =5087;
28007: waveform_sig_loopback =4068;
28008: waveform_sig_loopback =1416;
28009: waveform_sig_loopback =4218;
28010: waveform_sig_loopback =3276;
28011: waveform_sig_loopback =3096;
28012: waveform_sig_loopback =3742;
28013: waveform_sig_loopback =1853;
28014: waveform_sig_loopback =4601;
28015: waveform_sig_loopback =2584;
28016: waveform_sig_loopback =2430;
28017: waveform_sig_loopback =3728;
28018: waveform_sig_loopback =2762;
28019: waveform_sig_loopback =2397;
28020: waveform_sig_loopback =3157;
28021: waveform_sig_loopback =3503;
28022: waveform_sig_loopback =1566;
28023: waveform_sig_loopback =3243;
28024: waveform_sig_loopback =3064;
28025: waveform_sig_loopback =2248;
28026: waveform_sig_loopback =2191;
28027: waveform_sig_loopback =3483;
28028: waveform_sig_loopback =2351;
28029: waveform_sig_loopback =1272;
28030: waveform_sig_loopback =3555;
28031: waveform_sig_loopback =2911;
28032: waveform_sig_loopback =745;
28033: waveform_sig_loopback =2628;
28034: waveform_sig_loopback =3697;
28035: waveform_sig_loopback =1160;
28036: waveform_sig_loopback =1323;
28037: waveform_sig_loopback =3800;
28038: waveform_sig_loopback =1307;
28039: waveform_sig_loopback =2361;
28040: waveform_sig_loopback =3049;
28041: waveform_sig_loopback =-1710;
28042: waveform_sig_loopback =3857;
28043: waveform_sig_loopback =3086;
28044: waveform_sig_loopback =1150;
28045: waveform_sig_loopback =841;
28046: waveform_sig_loopback =987;
28047: waveform_sig_loopback =3651;
28048: waveform_sig_loopback =1840;
28049: waveform_sig_loopback =-102;
28050: waveform_sig_loopback =2475;
28051: waveform_sig_loopback =1135;
28052: waveform_sig_loopback =1828;
28053: waveform_sig_loopback =1435;
28054: waveform_sig_loopback =124;
28055: waveform_sig_loopback =3060;
28056: waveform_sig_loopback =333;
28057: waveform_sig_loopback =1055;
28058: waveform_sig_loopback =1677;
28059: waveform_sig_loopback =849;
28060: waveform_sig_loopback =925;
28061: waveform_sig_loopback =1131;
28062: waveform_sig_loopback =1633;
28063: waveform_sig_loopback =-152;
28064: waveform_sig_loopback =1422;
28065: waveform_sig_loopback =1190;
28066: waveform_sig_loopback =355;
28067: waveform_sig_loopback =335;
28068: waveform_sig_loopback =1686;
28069: waveform_sig_loopback =430;
28070: waveform_sig_loopback =-597;
28071: waveform_sig_loopback =1963;
28072: waveform_sig_loopback =769;
28073: waveform_sig_loopback =-1186;
28074: waveform_sig_loopback =1222;
28075: waveform_sig_loopback =1425;
28076: waveform_sig_loopback =-710;
28077: waveform_sig_loopback =-306;
28078: waveform_sig_loopback =1644;
28079: waveform_sig_loopback =-246;
28080: waveform_sig_loopback =389;
28081: waveform_sig_loopback =898;
28082: waveform_sig_loopback =-3158;
28083: waveform_sig_loopback =1718;
28084: waveform_sig_loopback =1375;
28085: waveform_sig_loopback =-734;
28086: waveform_sig_loopback =-1432;
28087: waveform_sig_loopback =-282;
28088: waveform_sig_loopback =1366;
28089: waveform_sig_loopback =-105;
28090: waveform_sig_loopback =-1632;
28091: waveform_sig_loopback =164;
28092: waveform_sig_loopback =-485;
28093: waveform_sig_loopback =-58;
28094: waveform_sig_loopback =-718;
28095: waveform_sig_loopback =-1332;
28096: waveform_sig_loopback =891;
28097: waveform_sig_loopback =-1578;
28098: waveform_sig_loopback =-599;
28099: waveform_sig_loopback =-516;
28100: waveform_sig_loopback =-890;
28101: waveform_sig_loopback =-930;
28102: waveform_sig_loopback =-858;
28103: waveform_sig_loopback =-215;
28104: waveform_sig_loopback =-1984;
28105: waveform_sig_loopback =-661;
28106: waveform_sig_loopback =-413;
28107: waveform_sig_loopback =-1748;
28108: waveform_sig_loopback =-1584;
28109: waveform_sig_loopback =220;
28110: waveform_sig_loopback =-2037;
28111: waveform_sig_loopback =-2091;
28112: waveform_sig_loopback =114;
28113: waveform_sig_loopback =-1516;
28114: waveform_sig_loopback =-2587;
28115: waveform_sig_loopback =-919;
28116: waveform_sig_loopback =-442;
28117: waveform_sig_loopback =-2441;
28118: waveform_sig_loopback =-2478;
28119: waveform_sig_loopback =35;
28120: waveform_sig_loopback =-2252;
28121: waveform_sig_loopback =-1579;
28122: waveform_sig_loopback =-898;
28123: waveform_sig_loopback =-5135;
28124: waveform_sig_loopback =-48;
28125: waveform_sig_loopback =-368;
28126: waveform_sig_loopback =-2969;
28127: waveform_sig_loopback =-3137;
28128: waveform_sig_loopback =-1934;
28129: waveform_sig_loopback =-819;
28130: waveform_sig_loopback =-1728;
28131: waveform_sig_loopback =-3633;
28132: waveform_sig_loopback =-1767;
28133: waveform_sig_loopback =-2077;
28134: waveform_sig_loopback =-2247;
28135: waveform_sig_loopback =-2478;
28136: waveform_sig_loopback =-2978;
28137: waveform_sig_loopback =-1299;
28138: waveform_sig_loopback =-3163;
28139: waveform_sig_loopback =-2507;
28140: waveform_sig_loopback =-2486;
28141: waveform_sig_loopback =-2465;
28142: waveform_sig_loopback =-3093;
28143: waveform_sig_loopback =-2523;
28144: waveform_sig_loopback =-1978;
28145: waveform_sig_loopback =-4080;
28146: waveform_sig_loopback =-2253;
28147: waveform_sig_loopback =-2273;
28148: waveform_sig_loopback =-3767;
28149: waveform_sig_loopback =-3067;
28150: waveform_sig_loopback =-1772;
28151: waveform_sig_loopback =-4004;
28152: waveform_sig_loopback =-3521;
28153: waveform_sig_loopback =-1973;
28154: waveform_sig_loopback =-3310;
28155: waveform_sig_loopback =-4229;
28156: waveform_sig_loopback =-2932;
28157: waveform_sig_loopback =-1996;
28158: waveform_sig_loopback =-4387;
28159: waveform_sig_loopback =-4348;
28160: waveform_sig_loopback =-1335;
28161: waveform_sig_loopback =-4521;
28162: waveform_sig_loopback =-3059;
28163: waveform_sig_loopback =-2638;
28164: waveform_sig_loopback =-7269;
28165: waveform_sig_loopback =-1216;
28166: waveform_sig_loopback =-2419;
28167: waveform_sig_loopback =-4940;
28168: waveform_sig_loopback =-4408;
28169: waveform_sig_loopback =-3990;
28170: waveform_sig_loopback =-2358;
28171: waveform_sig_loopback =-3401;
28172: waveform_sig_loopback =-5685;
28173: waveform_sig_loopback =-3006;
28174: waveform_sig_loopback =-3984;
28175: waveform_sig_loopback =-3952;
28176: waveform_sig_loopback =-3991;
28177: waveform_sig_loopback =-4860;
28178: waveform_sig_loopback =-2900;
28179: waveform_sig_loopback =-4738;
28180: waveform_sig_loopback =-4263;
28181: waveform_sig_loopback =-4076;
28182: waveform_sig_loopback =-4018;
28183: waveform_sig_loopback =-5025;
28184: waveform_sig_loopback =-3902;
28185: waveform_sig_loopback =-3695;
28186: waveform_sig_loopback =-5876;
28187: waveform_sig_loopback =-3433;
28188: waveform_sig_loopback =-4255;
28189: waveform_sig_loopback =-5327;
28190: waveform_sig_loopback =-4368;
28191: waveform_sig_loopback =-3812;
28192: waveform_sig_loopback =-5289;
28193: waveform_sig_loopback =-5085;
28194: waveform_sig_loopback =-3708;
28195: waveform_sig_loopback =-4613;
28196: waveform_sig_loopback =-6090;
28197: waveform_sig_loopback =-4348;
28198: waveform_sig_loopback =-3379;
28199: waveform_sig_loopback =-6404;
28200: waveform_sig_loopback =-5460;
28201: waveform_sig_loopback =-2889;
28202: waveform_sig_loopback =-6351;
28203: waveform_sig_loopback =-4023;
28204: waveform_sig_loopback =-4656;
28205: waveform_sig_loopback =-8667;
28206: waveform_sig_loopback =-2290;
28207: waveform_sig_loopback =-4405;
28208: waveform_sig_loopback =-6200;
28209: waveform_sig_loopback =-5857;
28210: waveform_sig_loopback =-5630;
28211: waveform_sig_loopback =-3420;
28212: waveform_sig_loopback =-5308;
28213: waveform_sig_loopback =-7077;
28214: waveform_sig_loopback =-4102;
28215: waveform_sig_loopback =-5894;
28216: waveform_sig_loopback =-5010;
28217: waveform_sig_loopback =-5534;
28218: waveform_sig_loopback =-6324;
28219: waveform_sig_loopback =-4099;
28220: waveform_sig_loopback =-6352;
28221: waveform_sig_loopback =-5598;
28222: waveform_sig_loopback =-5389;
28223: waveform_sig_loopback =-5398;
28224: waveform_sig_loopback =-6450;
28225: waveform_sig_loopback =-4963;
28226: waveform_sig_loopback =-5419;
28227: waveform_sig_loopback =-7169;
28228: waveform_sig_loopback =-4562;
28229: waveform_sig_loopback =-6078;
28230: waveform_sig_loopback =-6182;
28231: waveform_sig_loopback =-5883;
28232: waveform_sig_loopback =-5236;
28233: waveform_sig_loopback =-6181;
28234: waveform_sig_loopback =-6952;
28235: waveform_sig_loopback =-4555;
28236: waveform_sig_loopback =-5955;
28237: waveform_sig_loopback =-7689;
28238: waveform_sig_loopback =-4882;
28239: waveform_sig_loopback =-5155;
28240: waveform_sig_loopback =-7529;
28241: waveform_sig_loopback =-6378;
28242: waveform_sig_loopback =-4514;
28243: waveform_sig_loopback =-7307;
28244: waveform_sig_loopback =-5147;
28245: waveform_sig_loopback =-6188;
28246: waveform_sig_loopback =-9438;
28247: waveform_sig_loopback =-3453;
28248: waveform_sig_loopback =-5765;
28249: waveform_sig_loopback =-7125;
28250: waveform_sig_loopback =-7217;
28251: waveform_sig_loopback =-6675;
28252: waveform_sig_loopback =-4318;
28253: waveform_sig_loopback =-6729;
28254: waveform_sig_loopback =-7938;
28255: waveform_sig_loopback =-5133;
28256: waveform_sig_loopback =-7199;
28257: waveform_sig_loopback =-5706;
28258: waveform_sig_loopback =-6880;
28259: waveform_sig_loopback =-7309;
28260: waveform_sig_loopback =-4783;
28261: waveform_sig_loopback =-7820;
28262: waveform_sig_loopback =-6356;
28263: waveform_sig_loopback =-6298;
28264: waveform_sig_loopback =-6817;
28265: waveform_sig_loopback =-6965;
28266: waveform_sig_loopback =-6061;
28267: waveform_sig_loopback =-6563;
28268: waveform_sig_loopback =-7598;
28269: waveform_sig_loopback =-5918;
28270: waveform_sig_loopback =-6697;
28271: waveform_sig_loopback =-7112;
28272: waveform_sig_loopback =-7040;
28273: waveform_sig_loopback =-5674;
28274: waveform_sig_loopback =-7461;
28275: waveform_sig_loopback =-7684;
28276: waveform_sig_loopback =-5161;
28277: waveform_sig_loopback =-7254;
28278: waveform_sig_loopback =-8260;
28279: waveform_sig_loopback =-5679;
28280: waveform_sig_loopback =-6208;
28281: waveform_sig_loopback =-8143;
28282: waveform_sig_loopback =-7150;
28283: waveform_sig_loopback =-5366;
28284: waveform_sig_loopback =-8016;
28285: waveform_sig_loopback =-5882;
28286: waveform_sig_loopback =-7245;
28287: waveform_sig_loopback =-9815;
28288: waveform_sig_loopback =-4256;
28289: waveform_sig_loopback =-6566;
28290: waveform_sig_loopback =-7653;
28291: waveform_sig_loopback =-8217;
28292: waveform_sig_loopback =-6828;
28293: waveform_sig_loopback =-5155;
28294: waveform_sig_loopback =-7695;
28295: waveform_sig_loopback =-8078;
28296: waveform_sig_loopback =-6144;
28297: waveform_sig_loopback =-7607;
28298: waveform_sig_loopback =-6214;
28299: waveform_sig_loopback =-7877;
28300: waveform_sig_loopback =-7365;
28301: waveform_sig_loopback =-5676;
28302: waveform_sig_loopback =-8448;
28303: waveform_sig_loopback =-6462;
28304: waveform_sig_loopback =-7206;
28305: waveform_sig_loopback =-7150;
28306: waveform_sig_loopback =-7449;
28307: waveform_sig_loopback =-6754;
28308: waveform_sig_loopback =-6801;
28309: waveform_sig_loopback =-8229;
28310: waveform_sig_loopback =-6437;
28311: waveform_sig_loopback =-6875;
28312: waveform_sig_loopback =-7818;
28313: waveform_sig_loopback =-7277;
28314: waveform_sig_loopback =-6010;
28315: waveform_sig_loopback =-8121;
28316: waveform_sig_loopback =-7724;
28317: waveform_sig_loopback =-5610;
28318: waveform_sig_loopback =-7848;
28319: waveform_sig_loopback =-8302;
28320: waveform_sig_loopback =-6058;
28321: waveform_sig_loopback =-6730;
28322: waveform_sig_loopback =-8213;
28323: waveform_sig_loopback =-7546;
28324: waveform_sig_loopback =-5599;
28325: waveform_sig_loopback =-8234;
28326: waveform_sig_loopback =-6223;
28327: waveform_sig_loopback =-7418;
28328: waveform_sig_loopback =-10007;
28329: waveform_sig_loopback =-4680;
28330: waveform_sig_loopback =-6515;
28331: waveform_sig_loopback =-8187;
28332: waveform_sig_loopback =-8316;
28333: waveform_sig_loopback =-6789;
28334: waveform_sig_loopback =-5822;
28335: waveform_sig_loopback =-7468;
28336: waveform_sig_loopback =-8319;
28337: waveform_sig_loopback =-6534;
28338: waveform_sig_loopback =-7330;
28339: waveform_sig_loopback =-6715;
28340: waveform_sig_loopback =-7938;
28341: waveform_sig_loopback =-7231;
28342: waveform_sig_loopback =-6231;
28343: waveform_sig_loopback =-8139;
28344: waveform_sig_loopback =-6794;
28345: waveform_sig_loopback =-7557;
28346: waveform_sig_loopback =-6754;
28347: waveform_sig_loopback =-7731;
28348: waveform_sig_loopback =-6618;
28349: waveform_sig_loopback =-7091;
28350: waveform_sig_loopback =-8238;
28351: waveform_sig_loopback =-6065;
28352: waveform_sig_loopback =-6981;
28353: waveform_sig_loopback =-8060;
28354: waveform_sig_loopback =-6987;
28355: waveform_sig_loopback =-5790;
28356: waveform_sig_loopback =-8467;
28357: waveform_sig_loopback =-7329;
28358: waveform_sig_loopback =-5696;
28359: waveform_sig_loopback =-7800;
28360: waveform_sig_loopback =-7855;
28361: waveform_sig_loopback =-6453;
28362: waveform_sig_loopback =-6173;
28363: waveform_sig_loopback =-8206;
28364: waveform_sig_loopback =-7672;
28365: waveform_sig_loopback =-4956;
28366: waveform_sig_loopback =-8599;
28367: waveform_sig_loopback =-5656;
28368: waveform_sig_loopback =-7393;
28369: waveform_sig_loopback =-10154;
28370: waveform_sig_loopback =-3757;
28371: waveform_sig_loopback =-6674;
28372: waveform_sig_loopback =-8199;
28373: waveform_sig_loopback =-7597;
28374: waveform_sig_loopback =-6882;
28375: waveform_sig_loopback =-5325;
28376: waveform_sig_loopback =-7308;
28377: waveform_sig_loopback =-8240;
28378: waveform_sig_loopback =-5808;
28379: waveform_sig_loopback =-7264;
28380: waveform_sig_loopback =-6484;
28381: waveform_sig_loopback =-7349;
28382: waveform_sig_loopback =-6896;
28383: waveform_sig_loopback =-5906;
28384: waveform_sig_loopback =-7684;
28385: waveform_sig_loopback =-6475;
28386: waveform_sig_loopback =-6875;
28387: waveform_sig_loopback =-6352;
28388: waveform_sig_loopback =-7649;
28389: waveform_sig_loopback =-5851;
28390: waveform_sig_loopback =-6457;
28391: waveform_sig_loopback =-8103;
28392: waveform_sig_loopback =-5350;
28393: waveform_sig_loopback =-6808;
28394: waveform_sig_loopback =-7433;
28395: waveform_sig_loopback =-6073;
28396: waveform_sig_loopback =-6115;
28397: waveform_sig_loopback =-7393;
28398: waveform_sig_loopback =-6733;
28399: waveform_sig_loopback =-5432;
28400: waveform_sig_loopback =-6885;
28401: waveform_sig_loopback =-7679;
28402: waveform_sig_loopback =-5405;
28403: waveform_sig_loopback =-5636;
28404: waveform_sig_loopback =-8012;
28405: waveform_sig_loopback =-6456;
28406: waveform_sig_loopback =-4486;
28407: waveform_sig_loopback =-8122;
28408: waveform_sig_loopback =-4601;
28409: waveform_sig_loopback =-7136;
28410: waveform_sig_loopback =-9099;
28411: waveform_sig_loopback =-2932;
28412: waveform_sig_loopback =-6389;
28413: waveform_sig_loopback =-7073;
28414: waveform_sig_loopback =-6943;
28415: waveform_sig_loopback =-6213;
28416: waveform_sig_loopback =-4259;
28417: waveform_sig_loopback =-6789;
28418: waveform_sig_loopback =-7353;
28419: waveform_sig_loopback =-4921;
28420: waveform_sig_loopback =-6581;
28421: waveform_sig_loopback =-5490;
28422: waveform_sig_loopback =-6552;
28423: waveform_sig_loopback =-6168;
28424: waveform_sig_loopback =-4927;
28425: waveform_sig_loopback =-6732;
28426: waveform_sig_loopback =-5826;
28427: waveform_sig_loopback =-5703;
28428: waveform_sig_loopback =-5636;
28429: waveform_sig_loopback =-6832;
28430: waveform_sig_loopback =-4492;
28431: waveform_sig_loopback =-6206;
28432: waveform_sig_loopback =-6677;
28433: waveform_sig_loopback =-4365;
28434: waveform_sig_loopback =-6277;
28435: waveform_sig_loopback =-5909;
28436: waveform_sig_loopback =-5525;
28437: waveform_sig_loopback =-4937;
28438: waveform_sig_loopback =-6250;
28439: waveform_sig_loopback =-6106;
28440: waveform_sig_loopback =-4011;
28441: waveform_sig_loopback =-6105;
28442: waveform_sig_loopback =-6683;
28443: waveform_sig_loopback =-4063;
28444: waveform_sig_loopback =-4909;
28445: waveform_sig_loopback =-6858;
28446: waveform_sig_loopback =-5145;
28447: waveform_sig_loopback =-3701;
28448: waveform_sig_loopback =-6876;
28449: waveform_sig_loopback =-3329;
28450: waveform_sig_loopback =-6430;
28451: waveform_sig_loopback =-7572;
28452: waveform_sig_loopback =-1785;
28453: waveform_sig_loopback =-5473;
28454: waveform_sig_loopback =-5688;
28455: waveform_sig_loopback =-5955;
28456: waveform_sig_loopback =-4952;
28457: waveform_sig_loopback =-2834;
28458: waveform_sig_loopback =-5978;
28459: waveform_sig_loopback =-5884;
28460: waveform_sig_loopback =-3621;
28461: waveform_sig_loopback =-5712;
28462: waveform_sig_loopback =-3821;
28463: waveform_sig_loopback =-5631;
28464: waveform_sig_loopback =-4883;
28465: waveform_sig_loopback =-3358;
28466: waveform_sig_loopback =-5964;
28467: waveform_sig_loopback =-4213;
28468: waveform_sig_loopback =-4385;
28469: waveform_sig_loopback =-4765;
28470: waveform_sig_loopback =-4914;
28471: waveform_sig_loopback =-3544;
28472: waveform_sig_loopback =-4928;
28473: waveform_sig_loopback =-4924;
28474: waveform_sig_loopback =-3574;
28475: waveform_sig_loopback =-4476;
28476: waveform_sig_loopback =-4797;
28477: waveform_sig_loopback =-4162;
28478: waveform_sig_loopback =-3288;
28479: waveform_sig_loopback =-5245;
28480: waveform_sig_loopback =-4382;
28481: waveform_sig_loopback =-2626;
28482: waveform_sig_loopback =-4835;
28483: waveform_sig_loopback =-5151;
28484: waveform_sig_loopback =-2496;
28485: waveform_sig_loopback =-3614;
28486: waveform_sig_loopback =-5463;
28487: waveform_sig_loopback =-3379;
28488: waveform_sig_loopback =-2641;
28489: waveform_sig_loopback =-5112;
28490: waveform_sig_loopback =-1837;
28491: waveform_sig_loopback =-5426;
28492: waveform_sig_loopback =-5401;
28493: waveform_sig_loopback =-759;
28494: waveform_sig_loopback =-3815;
28495: waveform_sig_loopback =-4048;
28496: waveform_sig_loopback =-4872;
28497: waveform_sig_loopback =-2743;
28498: waveform_sig_loopback =-1719;
28499: waveform_sig_loopback =-4576;
28500: waveform_sig_loopback =-3888;
28501: waveform_sig_loopback =-2531;
28502: waveform_sig_loopback =-3800;
28503: waveform_sig_loopback =-2302;
28504: waveform_sig_loopback =-4356;
28505: waveform_sig_loopback =-2782;
28506: waveform_sig_loopback =-2125;
28507: waveform_sig_loopback =-4369;
28508: waveform_sig_loopback =-2273;
28509: waveform_sig_loopback =-3106;
28510: waveform_sig_loopback =-2921;
28511: waveform_sig_loopback =-3264;
28512: waveform_sig_loopback =-2071;
28513: waveform_sig_loopback =-3086;
28514: waveform_sig_loopback =-3301;
28515: waveform_sig_loopback =-2018;
28516: waveform_sig_loopback =-2602;
28517: waveform_sig_loopback =-3235;
28518: waveform_sig_loopback =-2411;
28519: waveform_sig_loopback =-1467;
28520: waveform_sig_loopback =-3892;
28521: waveform_sig_loopback =-2369;
28522: waveform_sig_loopback =-977;
28523: waveform_sig_loopback =-3432;
28524: waveform_sig_loopback =-3016;
28525: waveform_sig_loopback =-960;
28526: waveform_sig_loopback =-2007;
28527: waveform_sig_loopback =-3520;
28528: waveform_sig_loopback =-1766;
28529: waveform_sig_loopback =-913;
28530: waveform_sig_loopback =-3214;
28531: waveform_sig_loopback =-341;
28532: waveform_sig_loopback =-3621;
28533: waveform_sig_loopback =-3470;
28534: waveform_sig_loopback =769;
28535: waveform_sig_loopback =-1736;
28536: waveform_sig_loopback =-2738;
28537: waveform_sig_loopback =-2880;
28538: waveform_sig_loopback =-719;
28539: waveform_sig_loopback =-388;
28540: waveform_sig_loopback =-2414;
28541: waveform_sig_loopback =-2212;
28542: waveform_sig_loopback =-879;
28543: waveform_sig_loopback =-1642;
28544: waveform_sig_loopback =-849;
28545: waveform_sig_loopback =-2442;
28546: waveform_sig_loopback =-747;
28547: waveform_sig_loopback =-707;
28548: waveform_sig_loopback =-2218;
28549: waveform_sig_loopback =-609;
28550: waveform_sig_loopback =-1412;
28551: waveform_sig_loopback =-857;
28552: waveform_sig_loopback =-1673;
28553: waveform_sig_loopback =-127;
28554: waveform_sig_loopback =-1241;
28555: waveform_sig_loopback =-1609;
28556: waveform_sig_loopback =-26;
28557: waveform_sig_loopback =-766;
28558: waveform_sig_loopback =-1680;
28559: waveform_sig_loopback =-199;
28560: waveform_sig_loopback =197;
28561: waveform_sig_loopback =-2243;
28562: waveform_sig_loopback =-61;
28563: waveform_sig_loopback =479;
28564: waveform_sig_loopback =-1503;
28565: waveform_sig_loopback =-963;
28566: waveform_sig_loopback =617;
28567: waveform_sig_loopback =95;
28568: waveform_sig_loopback =-1834;
28569: waveform_sig_loopback =67;
28570: waveform_sig_loopback =1248;
28571: waveform_sig_loopback =-1720;
28572: waveform_sig_loopback =1773;
28573: waveform_sig_loopback =-1870;
28574: waveform_sig_loopback =-1681;
28575: waveform_sig_loopback =3021;
28576: waveform_sig_loopback =-114;
28577: waveform_sig_loopback =-1009;
28578: waveform_sig_loopback =-593;
28579: waveform_sig_loopback =918;
28580: waveform_sig_loopback =1520;
28581: waveform_sig_loopback =-443;
28582: waveform_sig_loopback =-528;
28583: waveform_sig_loopback =1273;
28584: waveform_sig_loopback =149;
28585: waveform_sig_loopback =840;
28586: waveform_sig_loopback =-214;
28587: waveform_sig_loopback =963;
28588: waveform_sig_loopback =1104;
28589: waveform_sig_loopback =-62;
28590: waveform_sig_loopback =1012;
28591: waveform_sig_loopback =669;
28592: waveform_sig_loopback =1021;
28593: waveform_sig_loopback =16;
28594: waveform_sig_loopback =2087;
28595: waveform_sig_loopback =403;
28596: waveform_sig_loopback =236;
28597: waveform_sig_loopback =2182;
28598: waveform_sig_loopback =754;
28599: waveform_sig_loopback =351;
28600: waveform_sig_loopback =1877;
28601: waveform_sig_loopback =1640;
28602: waveform_sig_loopback =11;
28603: waveform_sig_loopback =1770;
28604: waveform_sig_loopback =2212;
28605: waveform_sig_loopback =589;
28606: waveform_sig_loopback =737;
28607: waveform_sig_loopback =2601;
28608: waveform_sig_loopback =2006;
28609: waveform_sig_loopback =-182;
28610: waveform_sig_loopback =2283;
28611: waveform_sig_loopback =3046;
28612: waveform_sig_loopback =-77;
28613: waveform_sig_loopback =4049;
28614: waveform_sig_loopback =-375;
28615: waveform_sig_loopback =312;
28616: waveform_sig_loopback =5212;
28617: waveform_sig_loopback =1213;
28618: waveform_sig_loopback =1098;
28619: waveform_sig_loopback =1378;
28620: waveform_sig_loopback =2435;
28621: waveform_sig_loopback =3806;
28622: waveform_sig_loopback =987;
28623: waveform_sig_loopback =1418;
28624: waveform_sig_loopback =3391;
28625: waveform_sig_loopback =1583;
28626: waveform_sig_loopback =3012;
28627: waveform_sig_loopback =1509;
28628: waveform_sig_loopback =2699;
28629: waveform_sig_loopback =3165;
28630: waveform_sig_loopback =1605;
28631: waveform_sig_loopback =2894;
28632: waveform_sig_loopback =2651;
28633: waveform_sig_loopback =2626;
28634: waveform_sig_loopback =1966;
28635: waveform_sig_loopback =4012;
28636: waveform_sig_loopback =1994;
28637: waveform_sig_loopback =2284;
28638: waveform_sig_loopback =3990;
28639: waveform_sig_loopback =2319;
28640: waveform_sig_loopback =2471;
28641: waveform_sig_loopback =3702;
28642: waveform_sig_loopback =3229;
28643: waveform_sig_loopback =2109;
28644: waveform_sig_loopback =3339;
28645: waveform_sig_loopback =4141;
28646: waveform_sig_loopback =2421;
28647: waveform_sig_loopback =2233;
28648: waveform_sig_loopback =4832;
28649: waveform_sig_loopback =3509;
28650: waveform_sig_loopback =1465;
28651: waveform_sig_loopback =4583;
28652: waveform_sig_loopback =4211;
28653: waveform_sig_loopback =2016;
28654: waveform_sig_loopback =5960;
28655: waveform_sig_loopback =780;
28656: waveform_sig_loopback =2844;
28657: waveform_sig_loopback =6591;
28658: waveform_sig_loopback =2848;
28659: waveform_sig_loopback =3191;
28660: waveform_sig_loopback =2689;
28661: waveform_sig_loopback =4558;
28662: waveform_sig_loopback =5527;
28663: waveform_sig_loopback =2359;
28664: waveform_sig_loopback =3578;
28665: waveform_sig_loopback =4862;
28666: waveform_sig_loopback =3263;
28667: waveform_sig_loopback =4967;
28668: waveform_sig_loopback =2848;
28669: waveform_sig_loopback =4619;
28670: waveform_sig_loopback =4856;
28671: waveform_sig_loopback =3067;
28672: waveform_sig_loopback =4713;
28673: waveform_sig_loopback =4312;
28674: waveform_sig_loopback =4130;
28675: waveform_sig_loopback =3809;
28676: waveform_sig_loopback =5645;
28677: waveform_sig_loopback =3335;
28678: waveform_sig_loopback =4317;
28679: waveform_sig_loopback =5330;
28680: waveform_sig_loopback =3970;
28681: waveform_sig_loopback =4300;
28682: waveform_sig_loopback =4876;
28683: waveform_sig_loopback =5216;
28684: waveform_sig_loopback =3557;
28685: waveform_sig_loopback =4754;
28686: waveform_sig_loopback =6124;
28687: waveform_sig_loopback =3542;
28688: waveform_sig_loopback =3959;
28689: waveform_sig_loopback =6638;
28690: waveform_sig_loopback =4495;
28691: waveform_sig_loopback =3470;
28692: waveform_sig_loopback =5986;
28693: waveform_sig_loopback =5287;
28694: waveform_sig_loopback =4207;
28695: waveform_sig_loopback =7008;
28696: waveform_sig_loopback =2237;
28697: waveform_sig_loopback =4496;
28698: waveform_sig_loopback =7798;
28699: waveform_sig_loopback =4820;
28700: waveform_sig_loopback =4305;
28701: waveform_sig_loopback =4003;
28702: waveform_sig_loopback =6386;
28703: waveform_sig_loopback =6853;
28704: waveform_sig_loopback =3676;
28705: waveform_sig_loopback =5068;
28706: waveform_sig_loopback =6153;
28707: waveform_sig_loopback =4876;
28708: waveform_sig_loopback =6343;
28709: waveform_sig_loopback =3946;
28710: waveform_sig_loopback =6398;
28711: waveform_sig_loopback =6122;
28712: waveform_sig_loopback =4265;
28713: waveform_sig_loopback =6301;
28714: waveform_sig_loopback =5483;
28715: waveform_sig_loopback =5433;
28716: waveform_sig_loopback =5442;
28717: waveform_sig_loopback =6509;
28718: waveform_sig_loopback =4879;
28719: waveform_sig_loopback =5753;
28720: waveform_sig_loopback =6217;
28721: waveform_sig_loopback =5747;
28722: waveform_sig_loopback =5142;
28723: waveform_sig_loopback =6307;
28724: waveform_sig_loopback =6588;
28725: waveform_sig_loopback =4283;
28726: waveform_sig_loopback =6602;
28727: waveform_sig_loopback =7025;
28728: waveform_sig_loopback =4543;
28729: waveform_sig_loopback =5737;
28730: waveform_sig_loopback =7424;
28731: waveform_sig_loopback =5834;
28732: waveform_sig_loopback =4731;
28733: waveform_sig_loopback =7055;
28734: waveform_sig_loopback =6802;
28735: waveform_sig_loopback =5158;
28736: waveform_sig_loopback =8129;
28737: waveform_sig_loopback =3390;
28738: waveform_sig_loopback =5983;
28739: waveform_sig_loopback =8755;
28740: waveform_sig_loopback =5724;
28741: waveform_sig_loopback =5431;
28742: waveform_sig_loopback =5315;
28743: waveform_sig_loopback =7627;
28744: waveform_sig_loopback =7458;
28745: waveform_sig_loopback =4936;
28746: waveform_sig_loopback =6473;
28747: waveform_sig_loopback =6767;
28748: waveform_sig_loopback =6251;
28749: waveform_sig_loopback =7121;
28750: waveform_sig_loopback =5089;
28751: waveform_sig_loopback =7739;
28752: waveform_sig_loopback =6472;
28753: waveform_sig_loopback =5735;
28754: waveform_sig_loopback =7341;
28755: waveform_sig_loopback =6128;
28756: waveform_sig_loopback =6837;
28757: waveform_sig_loopback =6088;
28758: waveform_sig_loopback =7638;
28759: waveform_sig_loopback =5994;
28760: waveform_sig_loopback =6263;
28761: waveform_sig_loopback =7623;
28762: waveform_sig_loopback =6448;
28763: waveform_sig_loopback =5979;
28764: waveform_sig_loopback =7605;
28765: waveform_sig_loopback =7114;
28766: waveform_sig_loopback =5378;
28767: waveform_sig_loopback =7597;
28768: waveform_sig_loopback =7696;
28769: waveform_sig_loopback =5454;
28770: waveform_sig_loopback =6749;
28771: waveform_sig_loopback =8088;
28772: waveform_sig_loopback =6640;
28773: waveform_sig_loopback =5616;
28774: waveform_sig_loopback =7762;
28775: waveform_sig_loopback =7690;
28776: waveform_sig_loopback =5756;
28777: waveform_sig_loopback =8876;
28778: waveform_sig_loopback =4211;
28779: waveform_sig_loopback =6594;
28780: waveform_sig_loopback =9628;
28781: waveform_sig_loopback =6386;
28782: waveform_sig_loopback =5934;
28783: waveform_sig_loopback =6351;
28784: waveform_sig_loopback =8073;
28785: waveform_sig_loopback =8048;
28786: waveform_sig_loopback =5846;
28787: waveform_sig_loopback =6845;
28788: waveform_sig_loopback =7540;
28789: waveform_sig_loopback =6996;
28790: waveform_sig_loopback =7357;
28791: waveform_sig_loopback =6111;
28792: waveform_sig_loopback =8113;
28793: waveform_sig_loopback =6945;
28794: waveform_sig_loopback =6729;
28795: waveform_sig_loopback =7388;
28796: waveform_sig_loopback =7043;
28797: waveform_sig_loopback =7260;
28798: waveform_sig_loopback =6417;
28799: waveform_sig_loopback =8519;
28800: waveform_sig_loopback =6049;
28801: waveform_sig_loopback =6974;
28802: waveform_sig_loopback =8208;
28803: waveform_sig_loopback =6587;
28804: waveform_sig_loopback =6649;
28805: waveform_sig_loopback =8061;
28806: waveform_sig_loopback =7311;
28807: waveform_sig_loopback =5946;
28808: waveform_sig_loopback =8013;
28809: waveform_sig_loopback =7932;
28810: waveform_sig_loopback =5896;
28811: waveform_sig_loopback =7123;
28812: waveform_sig_loopback =8369;
28813: waveform_sig_loopback =7095;
28814: waveform_sig_loopback =5733;
28815: waveform_sig_loopback =8259;
28816: waveform_sig_loopback =8042;
28817: waveform_sig_loopback =5786;
28818: waveform_sig_loopback =9594;
28819: waveform_sig_loopback =4077;
28820: waveform_sig_loopback =7053;
28821: waveform_sig_loopback =10236;
28822: waveform_sig_loopback =5995;
28823: waveform_sig_loopback =6478;
28824: waveform_sig_loopback =6630;
28825: waveform_sig_loopback =8041;
28826: waveform_sig_loopback =8626;
28827: waveform_sig_loopback =5574;
28828: waveform_sig_loopback =7192;
28829: waveform_sig_loopback =7880;
28830: waveform_sig_loopback =6781;
28831: waveform_sig_loopback =7731;
28832: waveform_sig_loopback =6211;
28833: waveform_sig_loopback =8010;
28834: waveform_sig_loopback =7274;
28835: waveform_sig_loopback =6615;
28836: waveform_sig_loopback =7456;
28837: waveform_sig_loopback =7271;
28838: waveform_sig_loopback =7066;
28839: waveform_sig_loopback =6620;
28840: waveform_sig_loopback =8587;
28841: waveform_sig_loopback =5862;
28842: waveform_sig_loopback =7180;
28843: waveform_sig_loopback =8173;
28844: waveform_sig_loopback =6261;
28845: waveform_sig_loopback =6947;
28846: waveform_sig_loopback =7899;
28847: waveform_sig_loopback =7000;
28848: waveform_sig_loopback =6279;
28849: waveform_sig_loopback =7612;
28850: waveform_sig_loopback =7944;
28851: waveform_sig_loopback =5874;
28852: waveform_sig_loopback =6691;
28853: waveform_sig_loopback =8689;
28854: waveform_sig_loopback =6593;
28855: waveform_sig_loopback =5522;
28856: waveform_sig_loopback =8604;
28857: waveform_sig_loopback =7208;
28858: waveform_sig_loopback =6033;
28859: waveform_sig_loopback =9288;
28860: waveform_sig_loopback =3434;
28861: waveform_sig_loopback =7513;
28862: waveform_sig_loopback =9517;
28863: waveform_sig_loopback =5757;
28864: waveform_sig_loopback =6467;
28865: waveform_sig_loopback =6081;
28866: waveform_sig_loopback =8019;
28867: waveform_sig_loopback =8286;
28868: waveform_sig_loopback =5011;
28869: waveform_sig_loopback =7166;
28870: waveform_sig_loopback =7356;
28871: waveform_sig_loopback =6404;
28872: waveform_sig_loopback =7553;
28873: waveform_sig_loopback =5566;
28874: waveform_sig_loopback =7813;
28875: waveform_sig_loopback =6897;
28876: waveform_sig_loopback =6058;
28877: waveform_sig_loopback =7158;
28878: waveform_sig_loopback =6911;
28879: waveform_sig_loopback =6334;
28880: waveform_sig_loopback =6544;
28881: waveform_sig_loopback =7934;
28882: waveform_sig_loopback =5186;
28883: waveform_sig_loopback =7160;
28884: waveform_sig_loopback =7221;
28885: waveform_sig_loopback =5991;
28886: waveform_sig_loopback =6460;
28887: waveform_sig_loopback =7077;
28888: waveform_sig_loopback =6860;
28889: waveform_sig_loopback =5385;
28890: waveform_sig_loopback =7155;
28891: waveform_sig_loopback =7528;
28892: waveform_sig_loopback =4939;
28893: waveform_sig_loopback =6399;
28894: waveform_sig_loopback =8052;
28895: waveform_sig_loopback =5692;
28896: waveform_sig_loopback =5215;
28897: waveform_sig_loopback =7868;
28898: waveform_sig_loopback =6303;
28899: waveform_sig_loopback =5793;
28900: waveform_sig_loopback =8241;
28901: waveform_sig_loopback =2691;
28902: waveform_sig_loopback =7228;
28903: waveform_sig_loopback =8424;
28904: waveform_sig_loopback =5237;
28905: waveform_sig_loopback =5626;
28906: waveform_sig_loopback =5194;
28907: waveform_sig_loopback =7626;
28908: waveform_sig_loopback =7196;
28909: waveform_sig_loopback =4190;
28910: waveform_sig_loopback =6717;
28911: waveform_sig_loopback =6154;
28912: waveform_sig_loopback =5843;
28913: waveform_sig_loopback =6742;
28914: waveform_sig_loopback =4447;
28915: waveform_sig_loopback =7362;
28916: waveform_sig_loopback =5794;
28917: waveform_sig_loopback =5111;
28918: waveform_sig_loopback =6595;
28919: waveform_sig_loopback =5709;
28920: waveform_sig_loopback =5546;
28921: waveform_sig_loopback =5813;
28922: waveform_sig_loopback =6618;
28923: waveform_sig_loopback =4658;
28924: waveform_sig_loopback =6055;
28925: waveform_sig_loopback =6071;
28926: waveform_sig_loopback =5433;
28927: waveform_sig_loopback =5076;
28928: waveform_sig_loopback =6357;
28929: waveform_sig_loopback =5856;
28930: waveform_sig_loopback =4122;
28931: waveform_sig_loopback =6532;
28932: waveform_sig_loopback =6198;
28933: waveform_sig_loopback =3909;
28934: waveform_sig_loopback =5642;
28935: waveform_sig_loopback =6731;
28936: waveform_sig_loopback =4647;
28937: waveform_sig_loopback =4305;
28938: waveform_sig_loopback =6698;
28939: waveform_sig_loopback =5125;
28940: waveform_sig_loopback =4941;
28941: waveform_sig_loopback =6794;
28942: waveform_sig_loopback =1670;
28943: waveform_sig_loopback =6322;
28944: waveform_sig_loopback =6944;
28945: waveform_sig_loopback =4363;
28946: waveform_sig_loopback =4121;
28947: waveform_sig_loopback =4221;
28948: waveform_sig_loopback =6698;
28949: waveform_sig_loopback =5428;
28950: waveform_sig_loopback =3407;
28951: waveform_sig_loopback =5448;
28952: waveform_sig_loopback =4723;
28953: waveform_sig_loopback =5067;
28954: waveform_sig_loopback =4937;
28955: waveform_sig_loopback =3520;
28956: waveform_sig_loopback =6229;
28957: waveform_sig_loopback =4057;
28958: waveform_sig_loopback =4327;
28959: waveform_sig_loopback =4989;
28960: waveform_sig_loopback =4417;
28961: waveform_sig_loopback =4418;
28962: waveform_sig_loopback =4201;
28963: waveform_sig_loopback =5463;
28964: waveform_sig_loopback =3291;
28965: waveform_sig_loopback =4620;
28966: waveform_sig_loopback =4834;
28967: waveform_sig_loopback =3958;
28968: waveform_sig_loopback =3672;
28969: waveform_sig_loopback =5093;
28970: waveform_sig_loopback =4253;
28971: waveform_sig_loopback =2729;
28972: waveform_sig_loopback =5364;
28973: waveform_sig_loopback =4436;
28974: waveform_sig_loopback =2520;
28975: waveform_sig_loopback =4455;
28976: waveform_sig_loopback =4909;
28977: waveform_sig_loopback =3392;
28978: waveform_sig_loopback =2782;
28979: waveform_sig_loopback =5214;
28980: waveform_sig_loopback =3822;
28981: waveform_sig_loopback =3259;
28982: waveform_sig_loopback =5338;
28983: waveform_sig_loopback =247;
28984: waveform_sig_loopback =4788;
28985: waveform_sig_loopback =5649;
28986: waveform_sig_loopback =2625;
28987: waveform_sig_loopback =2490;
28988: waveform_sig_loopback =3107;
28989: waveform_sig_loopback =4917;
28990: waveform_sig_loopback =3941;
28991: waveform_sig_loopback =1982;
28992: waveform_sig_loopback =3631;
28993: waveform_sig_loopback =3479;
28994: waveform_sig_loopback =3392;
28995: waveform_sig_loopback =3237;
28996: waveform_sig_loopback =2306;
28997: waveform_sig_loopback =4376;
28998: waveform_sig_loopback =2566;
28999: waveform_sig_loopback =2900;
29000: waveform_sig_loopback =3169;
29001: waveform_sig_loopback =3090;
29002: waveform_sig_loopback =2672;
29003: waveform_sig_loopback =2599;
29004: waveform_sig_loopback =3981;
29005: waveform_sig_loopback =1537;
29006: waveform_sig_loopback =3033;
29007: waveform_sig_loopback =3364;
29008: waveform_sig_loopback =2144;
29009: waveform_sig_loopback =2158;
29010: waveform_sig_loopback =3656;
29011: waveform_sig_loopback =2222;
29012: waveform_sig_loopback =1452;
29013: waveform_sig_loopback =3678;
29014: waveform_sig_loopback =2541;
29015: waveform_sig_loopback =1209;
29016: waveform_sig_loopback =2583;
29017: waveform_sig_loopback =3378;
29018: waveform_sig_loopback =1723;
29019: waveform_sig_loopback =846;
29020: waveform_sig_loopback =3876;
29021: waveform_sig_loopback =1812;
29022: waveform_sig_loopback =1598;
29023: waveform_sig_loopback =3737;
29024: waveform_sig_loopback =-1749;
29025: waveform_sig_loopback =3325;
29026: waveform_sig_loopback =3860;
29027: waveform_sig_loopback =658;
29028: waveform_sig_loopback =949;
29029: waveform_sig_loopback =1399;
29030: waveform_sig_loopback =2948;
29031: waveform_sig_loopback =2384;
29032: waveform_sig_loopback =-31;
29033: waveform_sig_loopback =1999;
29034: waveform_sig_loopback =1832;
29035: waveform_sig_loopback =1334;
29036: waveform_sig_loopback =1628;
29037: waveform_sig_loopback =504;
29038: waveform_sig_loopback =2422;
29039: waveform_sig_loopback =884;
29040: waveform_sig_loopback =979;
29041: waveform_sig_loopback =1278;
29042: waveform_sig_loopback =1188;
29043: waveform_sig_loopback =806;
29044: waveform_sig_loopback =987;
29045: waveform_sig_loopback =2039;
29046: waveform_sig_loopback =-692;
29047: waveform_sig_loopback =1577;
29048: waveform_sig_loopback =1615;
29049: waveform_sig_loopback =-78;
29050: waveform_sig_loopback =536;
29051: waveform_sig_loopback =1690;
29052: waveform_sig_loopback =403;
29053: waveform_sig_loopback =-255;
29054: waveform_sig_loopback =1485;
29055: waveform_sig_loopback =905;
29056: waveform_sig_loopback =-672;
29057: waveform_sig_loopback =529;
29058: waveform_sig_loopback =1722;
29059: waveform_sig_loopback =-452;
29060: waveform_sig_loopback =-812;
29061: waveform_sig_loopback =2173;
29062: waveform_sig_loopback =-561;
29063: waveform_sig_loopback =244;
29064: waveform_sig_loopback =1619;
29065: waveform_sig_loopback =-3859;
29066: waveform_sig_loopback =1904;
29067: waveform_sig_loopback =1642;
29068: waveform_sig_loopback =-1207;
29069: waveform_sig_loopback =-857;
29070: waveform_sig_loopback =-681;
29071: waveform_sig_loopback =1260;
29072: waveform_sig_loopback =491;
29073: waveform_sig_loopback =-2241;
29074: waveform_sig_loopback =398;
29075: waveform_sig_loopback =-219;
29076: waveform_sig_loopback =-656;
29077: waveform_sig_loopback =-63;
29078: waveform_sig_loopback =-1696;
29079: waveform_sig_loopback =750;
29080: waveform_sig_loopback =-987;
29081: waveform_sig_loopback =-1238;
29082: waveform_sig_loopback =-219;
29083: waveform_sig_loopback =-696;
29084: waveform_sig_loopback =-1355;
29085: waveform_sig_loopback =-629;
29086: waveform_sig_loopback =-128;
29087: waveform_sig_loopback =-2262;
29088: waveform_sig_loopback =-336;
29089: waveform_sig_loopback =-697;
29090: waveform_sig_loopback =-1715;
29091: waveform_sig_loopback =-1203;
29092: waveform_sig_loopback =-377;
29093: waveform_sig_loopback =-1636;
29094: waveform_sig_loopback =-2048;
29095: waveform_sig_loopback =-398;
29096: waveform_sig_loopback =-902;
29097: waveform_sig_loopback =-2838;
29098: waveform_sig_loopback =-1243;
29099: waveform_sig_loopback =91;
29100: waveform_sig_loopback =-2844;
29101: waveform_sig_loopback =-2358;
29102: waveform_sig_loopback =272;
29103: waveform_sig_loopback =-2771;
29104: waveform_sig_loopback =-1098;
29105: waveform_sig_loopback =-908;
29106: waveform_sig_loopback =-5493;
29107: waveform_sig_loopback =451;
29108: waveform_sig_loopback =-845;
29109: waveform_sig_loopback =-2669;
29110: waveform_sig_loopback =-2889;
29111: waveform_sig_loopback =-2627;
29112: waveform_sig_loopback =-237;
29113: waveform_sig_loopback =-1919;
29114: waveform_sig_loopback =-3854;
29115: waveform_sig_loopback =-1291;
29116: waveform_sig_loopback =-2517;
29117: waveform_sig_loopback =-2028;
29118: waveform_sig_loopback =-2266;
29119: waveform_sig_loopback =-3496;
29120: waveform_sig_loopback =-878;
29121: waveform_sig_loopback =-3154;
29122: waveform_sig_loopback =-2777;
29123: waveform_sig_loopback =-2176;
29124: waveform_sig_loopback =-2567;
29125: waveform_sig_loopback =-3207;
29126: waveform_sig_loopback =-2245;
29127: waveform_sig_loopback =-2223;
29128: waveform_sig_loopback =-4037;
29129: waveform_sig_loopback =-1964;
29130: waveform_sig_loopback =-2812;
29131: waveform_sig_loopback =-3186;
29132: waveform_sig_loopback =-3300;
29133: waveform_sig_loopback =-2133;
29134: waveform_sig_loopback =-3171;
29135: waveform_sig_loopback =-4271;
29136: waveform_sig_loopback =-1799;
29137: waveform_sig_loopback =-2887;
29138: waveform_sig_loopback =-4821;
29139: waveform_sig_loopback =-2525;
29140: waveform_sig_loopback =-2144;
29141: waveform_sig_loopback =-4528;
29142: waveform_sig_loopback =-3869;
29143: waveform_sig_loopback =-1881;
29144: waveform_sig_loopback =-4254;
29145: waveform_sig_loopback =-2863;
29146: waveform_sig_loopback =-2967;
29147: waveform_sig_loopback =-6895;
29148: waveform_sig_loopback =-1475;
29149: waveform_sig_loopback =-2578;
29150: waveform_sig_loopback =-4329;
29151: waveform_sig_loopback =-4911;
29152: waveform_sig_loopback =-4034;
29153: waveform_sig_loopback =-2013;
29154: waveform_sig_loopback =-3794;
29155: waveform_sig_loopback =-5367;
29156: waveform_sig_loopback =-3096;
29157: waveform_sig_loopback =-4236;
29158: waveform_sig_loopback =-3597;
29159: waveform_sig_loopback =-4134;
29160: waveform_sig_loopback =-5066;
29161: waveform_sig_loopback =-2517;
29162: waveform_sig_loopback =-5039;
29163: waveform_sig_loopback =-4321;
29164: waveform_sig_loopback =-3795;
29165: waveform_sig_loopback =-4444;
29166: waveform_sig_loopback =-4649;
29167: waveform_sig_loopback =-3902;
29168: waveform_sig_loopback =-4120;
29169: waveform_sig_loopback =-5315;
29170: waveform_sig_loopback =-3918;
29171: waveform_sig_loopback =-4288;
29172: waveform_sig_loopback =-4723;
29173: waveform_sig_loopback =-5258;
29174: waveform_sig_loopback =-3246;
29175: waveform_sig_loopback =-5187;
29176: waveform_sig_loopback =-5790;
29177: waveform_sig_loopback =-2989;
29178: waveform_sig_loopback =-5070;
29179: waveform_sig_loopback =-5986;
29180: waveform_sig_loopback =-4063;
29181: waveform_sig_loopback =-3980;
29182: waveform_sig_loopback =-5760;
29183: waveform_sig_loopback =-5698;
29184: waveform_sig_loopback =-3204;
29185: waveform_sig_loopback =-5828;
29186: waveform_sig_loopback =-4495;
29187: waveform_sig_loopback =-4415;
29188: waveform_sig_loopback =-8453;
29189: waveform_sig_loopback =-2803;
29190: waveform_sig_loopback =-4103;
29191: waveform_sig_loopback =-5992;
29192: waveform_sig_loopback =-6295;
29193: waveform_sig_loopback =-5325;
29194: waveform_sig_loopback =-3533;
29195: waveform_sig_loopback =-5442;
29196: waveform_sig_loopback =-6599;
29197: waveform_sig_loopback =-4524;
29198: waveform_sig_loopback =-5735;
29199: waveform_sig_loopback =-4824;
29200: waveform_sig_loopback =-5847;
29201: waveform_sig_loopback =-6099;
29202: waveform_sig_loopback =-3981;
29203: waveform_sig_loopback =-6695;
29204: waveform_sig_loopback =-5209;
29205: waveform_sig_loopback =-5542;
29206: waveform_sig_loopback =-5689;
29207: waveform_sig_loopback =-5810;
29208: waveform_sig_loopback =-5724;
29209: waveform_sig_loopback =-4945;
29210: waveform_sig_loopback =-6954;
29211: waveform_sig_loopback =-5329;
29212: waveform_sig_loopback =-5163;
29213: waveform_sig_loopback =-6754;
29214: waveform_sig_loopback =-5991;
29215: waveform_sig_loopback =-4719;
29216: waveform_sig_loopback =-6856;
29217: waveform_sig_loopback =-6503;
29218: waveform_sig_loopback =-4702;
29219: waveform_sig_loopback =-6184;
29220: waveform_sig_loopback =-7299;
29221: waveform_sig_loopback =-5326;
29222: waveform_sig_loopback =-5101;
29223: waveform_sig_loopback =-7195;
29224: waveform_sig_loopback =-6750;
29225: waveform_sig_loopback =-4442;
29226: waveform_sig_loopback =-7058;
29227: waveform_sig_loopback =-5666;
29228: waveform_sig_loopback =-5724;
29229: waveform_sig_loopback =-9457;
29230: waveform_sig_loopback =-4062;
29231: waveform_sig_loopback =-5109;
29232: waveform_sig_loopback =-7298;
29233: waveform_sig_loopback =-7446;
29234: waveform_sig_loopback =-6170;
29235: waveform_sig_loopback =-4979;
29236: waveform_sig_loopback =-6276;
29237: waveform_sig_loopback =-7772;
29238: waveform_sig_loopback =-5854;
29239: waveform_sig_loopback =-6362;
29240: waveform_sig_loopback =-6247;
29241: waveform_sig_loopback =-6902;
29242: waveform_sig_loopback =-6845;
29243: waveform_sig_loopback =-5478;
29244: waveform_sig_loopback =-7342;
29245: waveform_sig_loopback =-6358;
29246: waveform_sig_loopback =-6755;
29247: waveform_sig_loopback =-6203;
29248: waveform_sig_loopback =-7291;
29249: waveform_sig_loopback =-6289;
29250: waveform_sig_loopback =-5958;
29251: waveform_sig_loopback =-8219;
29252: waveform_sig_loopback =-5702;
29253: waveform_sig_loopback =-6460;
29254: waveform_sig_loopback =-7622;
29255: waveform_sig_loopback =-6604;
29256: waveform_sig_loopback =-5832;
29257: waveform_sig_loopback =-7589;
29258: waveform_sig_loopback =-7312;
29259: waveform_sig_loopback =-5595;
29260: waveform_sig_loopback =-7005;
29261: waveform_sig_loopback =-8073;
29262: waveform_sig_loopback =-6146;
29263: waveform_sig_loopback =-5872;
29264: waveform_sig_loopback =-8015;
29265: waveform_sig_loopback =-7620;
29266: waveform_sig_loopback =-4957;
29267: waveform_sig_loopback =-8009;
29268: waveform_sig_loopback =-6301;
29269: waveform_sig_loopback =-6413;
29270: waveform_sig_loopback =-10460;
29271: waveform_sig_loopback =-4381;
29272: waveform_sig_loopback =-5948;
29273: waveform_sig_loopback =-8387;
29274: waveform_sig_loopback =-7609;
29275: waveform_sig_loopback =-7212;
29276: waveform_sig_loopback =-5591;
29277: waveform_sig_loopback =-6729;
29278: waveform_sig_loopback =-8951;
29279: waveform_sig_loopback =-5972;
29280: waveform_sig_loopback =-7290;
29281: waveform_sig_loopback =-6976;
29282: waveform_sig_loopback =-7123;
29283: waveform_sig_loopback =-7799;
29284: waveform_sig_loopback =-5905;
29285: waveform_sig_loopback =-7807;
29286: waveform_sig_loopback =-7182;
29287: waveform_sig_loopback =-6929;
29288: waveform_sig_loopback =-6938;
29289: waveform_sig_loopback =-7854;
29290: waveform_sig_loopback =-6423;
29291: waveform_sig_loopback =-6824;
29292: waveform_sig_loopback =-8457;
29293: waveform_sig_loopback =-6085;
29294: waveform_sig_loopback =-7041;
29295: waveform_sig_loopback =-7953;
29296: waveform_sig_loopback =-6910;
29297: waveform_sig_loopback =-6356;
29298: waveform_sig_loopback =-7989;
29299: waveform_sig_loopback =-7532;
29300: waveform_sig_loopback =-6177;
29301: waveform_sig_loopback =-7226;
29302: waveform_sig_loopback =-8513;
29303: waveform_sig_loopback =-6511;
29304: waveform_sig_loopback =-5989;
29305: waveform_sig_loopback =-8824;
29306: waveform_sig_loopback =-7581;
29307: waveform_sig_loopback =-5287;
29308: waveform_sig_loopback =-8821;
29309: waveform_sig_loopback =-5900;
29310: waveform_sig_loopback =-7397;
29311: waveform_sig_loopback =-10572;
29312: waveform_sig_loopback =-4095;
29313: waveform_sig_loopback =-6954;
29314: waveform_sig_loopback =-8163;
29315: waveform_sig_loopback =-7951;
29316: waveform_sig_loopback =-7582;
29317: waveform_sig_loopback =-5169;
29318: waveform_sig_loopback =-7571;
29319: waveform_sig_loopback =-8784;
29320: waveform_sig_loopback =-5892;
29321: waveform_sig_loopback =-7844;
29322: waveform_sig_loopback =-6587;
29323: waveform_sig_loopback =-7533;
29324: waveform_sig_loopback =-7846;
29325: waveform_sig_loopback =-5732;
29326: waveform_sig_loopback =-8194;
29327: waveform_sig_loopback =-7068;
29328: waveform_sig_loopback =-6958;
29329: waveform_sig_loopback =-7073;
29330: waveform_sig_loopback =-7906;
29331: waveform_sig_loopback =-6323;
29332: waveform_sig_loopback =-7064;
29333: waveform_sig_loopback =-8260;
29334: waveform_sig_loopback =-6003;
29335: waveform_sig_loopback =-7420;
29336: waveform_sig_loopback =-7523;
29337: waveform_sig_loopback =-7024;
29338: waveform_sig_loopback =-6442;
29339: waveform_sig_loopback =-7629;
29340: waveform_sig_loopback =-7912;
29341: waveform_sig_loopback =-5632;
29342: waveform_sig_loopback =-7322;
29343: waveform_sig_loopback =-8642;
29344: waveform_sig_loopback =-5794;
29345: waveform_sig_loopback =-6336;
29346: waveform_sig_loopback =-8526;
29347: waveform_sig_loopback =-7098;
29348: waveform_sig_loopback =-5439;
29349: waveform_sig_loopback =-8396;
29350: waveform_sig_loopback =-5544;
29351: waveform_sig_loopback =-7570;
29352: waveform_sig_loopback =-9838;
29353: waveform_sig_loopback =-3934;
29354: waveform_sig_loopback =-6902;
29355: waveform_sig_loopback =-7505;
29356: waveform_sig_loopback =-8007;
29357: waveform_sig_loopback =-6950;
29358: waveform_sig_loopback =-4808;
29359: waveform_sig_loopback =-7698;
29360: waveform_sig_loopback =-7971;
29361: waveform_sig_loopback =-5767;
29362: waveform_sig_loopback =-7564;
29363: waveform_sig_loopback =-5929;
29364: waveform_sig_loopback =-7592;
29365: waveform_sig_loopback =-7139;
29366: waveform_sig_loopback =-5370;
29367: waveform_sig_loopback =-8026;
29368: waveform_sig_loopback =-6383;
29369: waveform_sig_loopback =-6684;
29370: waveform_sig_loopback =-6737;
29371: waveform_sig_loopback =-7253;
29372: waveform_sig_loopback =-5889;
29373: waveform_sig_loopback =-6784;
29374: waveform_sig_loopback =-7542;
29375: waveform_sig_loopback =-5684;
29376: waveform_sig_loopback =-6819;
29377: waveform_sig_loopback =-6909;
29378: waveform_sig_loopback =-6800;
29379: waveform_sig_loopback =-5527;
29380: waveform_sig_loopback =-7358;
29381: waveform_sig_loopback =-7308;
29382: waveform_sig_loopback =-4739;
29383: waveform_sig_loopback =-7212;
29384: waveform_sig_loopback =-7690;
29385: waveform_sig_loopback =-5071;
29386: waveform_sig_loopback =-6099;
29387: waveform_sig_loopback =-7586;
29388: waveform_sig_loopback =-6529;
29389: waveform_sig_loopback =-4864;
29390: waveform_sig_loopback =-7586;
29391: waveform_sig_loopback =-5217;
29392: waveform_sig_loopback =-6801;
29393: waveform_sig_loopback =-8867;
29394: waveform_sig_loopback =-3527;
29395: waveform_sig_loopback =-6111;
29396: waveform_sig_loopback =-6835;
29397: waveform_sig_loopback =-7223;
29398: waveform_sig_loopback =-5943;
29399: waveform_sig_loopback =-4482;
29400: waveform_sig_loopback =-6826;
29401: waveform_sig_loopback =-6881;
29402: waveform_sig_loopback =-5377;
29403: waveform_sig_loopback =-6606;
29404: waveform_sig_loopback =-5120;
29405: waveform_sig_loopback =-6910;
29406: waveform_sig_loopback =-5995;
29407: waveform_sig_loopback =-4906;
29408: waveform_sig_loopback =-7064;
29409: waveform_sig_loopback =-5268;
29410: waveform_sig_loopback =-6100;
29411: waveform_sig_loopback =-5786;
29412: waveform_sig_loopback =-6227;
29413: waveform_sig_loopback =-5136;
29414: waveform_sig_loopback =-5747;
29415: waveform_sig_loopback =-6698;
29416: waveform_sig_loopback =-4847;
29417: waveform_sig_loopback =-5537;
29418: waveform_sig_loopback =-6368;
29419: waveform_sig_loopback =-5601;
29420: waveform_sig_loopback =-4405;
29421: waveform_sig_loopback =-6710;
29422: waveform_sig_loopback =-5916;
29423: waveform_sig_loopback =-3858;
29424: waveform_sig_loopback =-6342;
29425: waveform_sig_loopback =-6283;
29426: waveform_sig_loopback =-4308;
29427: waveform_sig_loopback =-5001;
29428: waveform_sig_loopback =-6335;
29429: waveform_sig_loopback =-5665;
29430: waveform_sig_loopback =-3589;
29431: waveform_sig_loopback =-6484;
29432: waveform_sig_loopback =-4022;
29433: waveform_sig_loopback =-5710;
29434: waveform_sig_loopback =-7878;
29435: waveform_sig_loopback =-2225;
29436: waveform_sig_loopback =-4668;
29437: waveform_sig_loopback =-6222;
29438: waveform_sig_loopback =-5872;
29439: waveform_sig_loopback =-4656;
29440: waveform_sig_loopback =-3466;
29441: waveform_sig_loopback =-5368;
29442: waveform_sig_loopback =-6060;
29443: waveform_sig_loopback =-3966;
29444: waveform_sig_loopback =-5190;
29445: waveform_sig_loopback =-4190;
29446: waveform_sig_loopback =-5566;
29447: waveform_sig_loopback =-4596;
29448: waveform_sig_loopback =-3762;
29449: waveform_sig_loopback =-5715;
29450: waveform_sig_loopback =-4043;
29451: waveform_sig_loopback =-4841;
29452: waveform_sig_loopback =-4219;
29453: waveform_sig_loopback =-5120;
29454: waveform_sig_loopback =-3799;
29455: waveform_sig_loopback =-4212;
29456: waveform_sig_loopback =-5541;
29457: waveform_sig_loopback =-3301;
29458: waveform_sig_loopback =-4156;
29459: waveform_sig_loopback =-5339;
29460: waveform_sig_loopback =-3697;
29461: waveform_sig_loopback =-3425;
29462: waveform_sig_loopback =-5387;
29463: waveform_sig_loopback =-4014;
29464: waveform_sig_loopback =-3000;
29465: waveform_sig_loopback =-4687;
29466: waveform_sig_loopback =-4968;
29467: waveform_sig_loopback =-3015;
29468: waveform_sig_loopback =-3233;
29469: waveform_sig_loopback =-5327;
29470: waveform_sig_loopback =-3943;
29471: waveform_sig_loopback =-2023;
29472: waveform_sig_loopback =-5403;
29473: waveform_sig_loopback =-2127;
29474: waveform_sig_loopback =-4643;
29475: waveform_sig_loopback =-6231;
29476: waveform_sig_loopback =-421;
29477: waveform_sig_loopback =-3579;
29478: waveform_sig_loopback =-4654;
29479: waveform_sig_loopback =-4209;
29480: waveform_sig_loopback =-3177;
29481: waveform_sig_loopback =-1856;
29482: waveform_sig_loopback =-3917;
29483: waveform_sig_loopback =-4495;
29484: waveform_sig_loopback =-2265;
29485: waveform_sig_loopback =-3607;
29486: waveform_sig_loopback =-2793;
29487: waveform_sig_loopback =-3735;
29488: waveform_sig_loopback =-3090;
29489: waveform_sig_loopback =-2298;
29490: waveform_sig_loopback =-3798;
29491: waveform_sig_loopback =-2810;
29492: waveform_sig_loopback =-2933;
29493: waveform_sig_loopback =-2598;
29494: waveform_sig_loopback =-3846;
29495: waveform_sig_loopback =-1651;
29496: waveform_sig_loopback =-3036;
29497: waveform_sig_loopback =-3831;
29498: waveform_sig_loopback =-1397;
29499: waveform_sig_loopback =-2983;
29500: waveform_sig_loopback =-3203;
29501: waveform_sig_loopback =-2137;
29502: waveform_sig_loopback =-2020;
29503: waveform_sig_loopback =-3348;
29504: waveform_sig_loopback =-2590;
29505: waveform_sig_loopback =-1294;
29506: waveform_sig_loopback =-2881;
29507: waveform_sig_loopback =-3412;
29508: waveform_sig_loopback =-1092;
29509: waveform_sig_loopback =-1616;
29510: waveform_sig_loopback =-3805;
29511: waveform_sig_loopback =-1835;
29512: waveform_sig_loopback =-545;
29513: waveform_sig_loopback =-3762;
29514: waveform_sig_loopback =28;
29515: waveform_sig_loopback =-3455;
29516: waveform_sig_loopback =-4124;
29517: waveform_sig_loopback =1486;
29518: waveform_sig_loopback =-2235;
29519: waveform_sig_loopback =-2593;
29520: waveform_sig_loopback =-2522;
29521: waveform_sig_loopback =-1489;
29522: waveform_sig_loopback =183;
29523: waveform_sig_loopback =-2473;
29524: waveform_sig_loopback =-2618;
29525: waveform_sig_loopback =-297;
29526: waveform_sig_loopback =-2117;
29527: waveform_sig_loopback =-745;
29528: waveform_sig_loopback =-2000;
29529: waveform_sig_loopback =-1460;
29530: waveform_sig_loopback =-177;
29531: waveform_sig_loopback =-2194;
29532: waveform_sig_loopback =-1070;
29533: waveform_sig_loopback =-811;
29534: waveform_sig_loopback =-1199;
29535: waveform_sig_loopback =-1761;
29536: waveform_sig_loopback =263;
29537: waveform_sig_loopback =-1632;
29538: waveform_sig_loopback =-1422;
29539: waveform_sig_loopback =80;
29540: waveform_sig_loopback =-1149;
29541: waveform_sig_loopback =-1093;
29542: waveform_sig_loopback =-622;
29543: waveform_sig_loopback =134;
29544: waveform_sig_loopback =-1639;
29545: waveform_sig_loopback =-715;
29546: waveform_sig_loopback =742;
29547: waveform_sig_loopback =-1276;
29548: waveform_sig_loopback =-1412;
29549: waveform_sig_loopback =860;
29550: waveform_sig_loopback =101;
29551: waveform_sig_loopback =-2010;
29552: waveform_sig_loopback =346;
29553: waveform_sig_loopback =1044;
29554: waveform_sig_loopback =-1837;
29555: waveform_sig_loopback =2185;
29556: waveform_sig_loopback =-2218;
29557: waveform_sig_loopback =-1678;
29558: waveform_sig_loopback =3201;
29559: waveform_sig_loopback =-622;
29560: waveform_sig_loopback =-321;
29561: waveform_sig_loopback =-1103;
29562: waveform_sig_loopback =762;
29563: waveform_sig_loopback =2117;
29564: waveform_sig_loopback =-1130;
29565: waveform_sig_loopback =-127;
29566: waveform_sig_loopback =1226;
29567: waveform_sig_loopback =-277;
29568: waveform_sig_loopback =1450;
29569: waveform_sig_loopback =-674;
29570: waveform_sig_loopback =877;
29571: waveform_sig_loopback =1596;
29572: waveform_sig_loopback =-564;
29573: waveform_sig_loopback =1232;
29574: waveform_sig_loopback =789;
29575: waveform_sig_loopback =756;
29576: waveform_sig_loopback =306;
29577: waveform_sig_loopback =1923;
29578: waveform_sig_loopback =330;
29579: waveform_sig_loopback =552;
29580: waveform_sig_loopback =1822;
29581: waveform_sig_loopback =819;
29582: waveform_sig_loopback =744;
29583: waveform_sig_loopback =1260;
29584: waveform_sig_loopback =2051;
29585: waveform_sig_loopback =141;
29586: waveform_sig_loopback =1182;
29587: waveform_sig_loopback =2800;
29588: waveform_sig_loopback =335;
29589: waveform_sig_loopback =586;
29590: waveform_sig_loopback =2999;
29591: waveform_sig_loopback =1473;
29592: waveform_sig_loopback =202;
29593: waveform_sig_loopback =2240;
29594: waveform_sig_loopback =2593;
29595: waveform_sig_loopback =542;
29596: waveform_sig_loopback =3668;
29597: waveform_sig_loopback =-317;
29598: waveform_sig_loopback =586;
29599: waveform_sig_loopback =4649;
29600: waveform_sig_loopback =1714;
29601: waveform_sig_loopback =1211;
29602: waveform_sig_loopback =768;
29603: waveform_sig_loopback =3050;
29604: waveform_sig_loopback =3521;
29605: waveform_sig_loopback =931;
29606: waveform_sig_loopback =1766;
29607: waveform_sig_loopback =2855;
29608: waveform_sig_loopback =1924;
29609: waveform_sig_loopback =3146;
29610: waveform_sig_loopback =1105;
29611: waveform_sig_loopback =2981;
29612: waveform_sig_loopback =3141;
29613: waveform_sig_loopback =1415;
29614: waveform_sig_loopback =3117;
29615: waveform_sig_loopback =2442;
29616: waveform_sig_loopback =2632;
29617: waveform_sig_loopback =2204;
29618: waveform_sig_loopback =3625;
29619: waveform_sig_loopback =2184;
29620: waveform_sig_loopback =2438;
29621: waveform_sig_loopback =3439;
29622: waveform_sig_loopback =2934;
29623: waveform_sig_loopback =2215;
29624: waveform_sig_loopback =3242;
29625: waveform_sig_loopback =4038;
29626: waveform_sig_loopback =1475;
29627: waveform_sig_loopback =3491;
29628: waveform_sig_loopback =4331;
29629: waveform_sig_loopback =1973;
29630: waveform_sig_loopback =2776;
29631: waveform_sig_loopback =4390;
29632: waveform_sig_loopback =3442;
29633: waveform_sig_loopback =2023;
29634: waveform_sig_loopback =3871;
29635: waveform_sig_loopback =4580;
29636: waveform_sig_loopback =2139;
29637: waveform_sig_loopback =5392;
29638: waveform_sig_loopback =1504;
29639: waveform_sig_loopback =2231;
29640: waveform_sig_loopback =6525;
29641: waveform_sig_loopback =3404;
29642: waveform_sig_loopback =2637;
29643: waveform_sig_loopback =2909;
29644: waveform_sig_loopback =4582;
29645: waveform_sig_loopback =5139;
29646: waveform_sig_loopback =2799;
29647: waveform_sig_loopback =3356;
29648: waveform_sig_loopback =4672;
29649: waveform_sig_loopback =3595;
29650: waveform_sig_loopback =4710;
29651: waveform_sig_loopback =2886;
29652: waveform_sig_loopback =4738;
29653: waveform_sig_loopback =4615;
29654: waveform_sig_loopback =3177;
29655: waveform_sig_loopback =4827;
29656: waveform_sig_loopback =3944;
29657: waveform_sig_loopback =4471;
29658: waveform_sig_loopback =3714;
29659: waveform_sig_loopback =5233;
29660: waveform_sig_loopback =4067;
29661: waveform_sig_loopback =3686;
29662: waveform_sig_loopback =5358;
29663: waveform_sig_loopback =4487;
29664: waveform_sig_loopback =3502;
29665: waveform_sig_loopback =5389;
29666: waveform_sig_loopback =5048;
29667: waveform_sig_loopback =3256;
29668: waveform_sig_loopback =5314;
29669: waveform_sig_loopback =5441;
29670: waveform_sig_loopback =3950;
29671: waveform_sig_loopback =4110;
29672: waveform_sig_loopback =6018;
29673: waveform_sig_loopback =5111;
29674: waveform_sig_loopback =3234;
29675: waveform_sig_loopback =5735;
29676: waveform_sig_loopback =5924;
29677: waveform_sig_loopback =3606;
29678: waveform_sig_loopback =7109;
29679: waveform_sig_loopback =2650;
29680: waveform_sig_loopback =4017;
29681: waveform_sig_loopback =8019;
29682: waveform_sig_loopback =4742;
29683: waveform_sig_loopback =4095;
29684: waveform_sig_loopback =4434;
29685: waveform_sig_loopback =6146;
29686: waveform_sig_loopback =6549;
29687: waveform_sig_loopback =4260;
29688: waveform_sig_loopback =4691;
29689: waveform_sig_loopback =6158;
29690: waveform_sig_loopback =5191;
29691: waveform_sig_loopback =5754;
29692: waveform_sig_loopback =4603;
29693: waveform_sig_loopback =6090;
29694: waveform_sig_loopback =5845;
29695: waveform_sig_loopback =4951;
29696: waveform_sig_loopback =5785;
29697: waveform_sig_loopback =5660;
29698: waveform_sig_loopback =5762;
29699: waveform_sig_loopback =4783;
29700: waveform_sig_loopback =7134;
29701: waveform_sig_loopback =4796;
29702: waveform_sig_loopback =5344;
29703: waveform_sig_loopback =6844;
29704: waveform_sig_loopback =5284;
29705: waveform_sig_loopback =5309;
29706: waveform_sig_loopback =6497;
29707: waveform_sig_loopback =6263;
29708: waveform_sig_loopback =4703;
29709: waveform_sig_loopback =6441;
29710: waveform_sig_loopback =6828;
29711: waveform_sig_loopback =5043;
29712: waveform_sig_loopback =5417;
29713: waveform_sig_loopback =7277;
29714: waveform_sig_loopback =6240;
29715: waveform_sig_loopback =4356;
29716: waveform_sig_loopback =7085;
29717: waveform_sig_loopback =7065;
29718: waveform_sig_loopback =4604;
29719: waveform_sig_loopback =8487;
29720: waveform_sig_loopback =3485;
29721: waveform_sig_loopback =5413;
29722: waveform_sig_loopback =9311;
29723: waveform_sig_loopback =5440;
29724: waveform_sig_loopback =5464;
29725: waveform_sig_loopback =5634;
29726: waveform_sig_loopback =6970;
29727: waveform_sig_loopback =7914;
29728: waveform_sig_loopback =5036;
29729: waveform_sig_loopback =5871;
29730: waveform_sig_loopback =7480;
29731: waveform_sig_loopback =5817;
29732: waveform_sig_loopback =7153;
29733: waveform_sig_loopback =5571;
29734: waveform_sig_loopback =6857;
29735: waveform_sig_loopback =7244;
29736: waveform_sig_loopback =5636;
29737: waveform_sig_loopback =6907;
29738: waveform_sig_loopback =6590;
29739: waveform_sig_loopback =6422;
29740: waveform_sig_loopback =6274;
29741: waveform_sig_loopback =7894;
29742: waveform_sig_loopback =5367;
29743: waveform_sig_loopback =6525;
29744: waveform_sig_loopback =7862;
29745: waveform_sig_loopback =6148;
29746: waveform_sig_loopback =6180;
29747: waveform_sig_loopback =7314;
29748: waveform_sig_loopback =7271;
29749: waveform_sig_loopback =5646;
29750: waveform_sig_loopback =7072;
29751: waveform_sig_loopback =7790;
29752: waveform_sig_loopback =5890;
29753: waveform_sig_loopback =6184;
29754: waveform_sig_loopback =8239;
29755: waveform_sig_loopback =6882;
29756: waveform_sig_loopback =5207;
29757: waveform_sig_loopback =8193;
29758: waveform_sig_loopback =7390;
29759: waveform_sig_loopback =5626;
29760: waveform_sig_loopback =9488;
29761: waveform_sig_loopback =3639;
29762: waveform_sig_loopback =6723;
29763: waveform_sig_loopback =9841;
29764: waveform_sig_loopback =5959;
29765: waveform_sig_loopback =6485;
29766: waveform_sig_loopback =5909;
29767: waveform_sig_loopback =7990;
29768: waveform_sig_loopback =8653;
29769: waveform_sig_loopback =5202;
29770: waveform_sig_loopback =7043;
29771: waveform_sig_loopback =7777;
29772: waveform_sig_loopback =6433;
29773: waveform_sig_loopback =7979;
29774: waveform_sig_loopback =5713;
29775: waveform_sig_loopback =7933;
29776: waveform_sig_loopback =7583;
29777: waveform_sig_loopback =6013;
29778: waveform_sig_loopback =7705;
29779: waveform_sig_loopback =7134;
29780: waveform_sig_loopback =6900;
29781: waveform_sig_loopback =6770;
29782: waveform_sig_loopback =8321;
29783: waveform_sig_loopback =6040;
29784: waveform_sig_loopback =7224;
29785: waveform_sig_loopback =7910;
29786: waveform_sig_loopback =6614;
29787: waveform_sig_loopback =6944;
29788: waveform_sig_loopback =7598;
29789: waveform_sig_loopback =7614;
29790: waveform_sig_loopback =6015;
29791: waveform_sig_loopback =7513;
29792: waveform_sig_loopback =8486;
29793: waveform_sig_loopback =5737;
29794: waveform_sig_loopback =6757;
29795: waveform_sig_loopback =8941;
29796: waveform_sig_loopback =6609;
29797: waveform_sig_loopback =5942;
29798: waveform_sig_loopback =8447;
29799: waveform_sig_loopback =7497;
29800: waveform_sig_loopback =6388;
29801: waveform_sig_loopback =9174;
29802: waveform_sig_loopback =4101;
29803: waveform_sig_loopback =7329;
29804: waveform_sig_loopback =9643;
29805: waveform_sig_loopback =6507;
29806: waveform_sig_loopback =6540;
29807: waveform_sig_loopback =6120;
29808: waveform_sig_loopback =8504;
29809: waveform_sig_loopback =8491;
29810: waveform_sig_loopback =5442;
29811: waveform_sig_loopback =7476;
29812: waveform_sig_loopback =7553;
29813: waveform_sig_loopback =6835;
29814: waveform_sig_loopback =8085;
29815: waveform_sig_loopback =5587;
29816: waveform_sig_loopback =8468;
29817: waveform_sig_loopback =7275;
29818: waveform_sig_loopback =6233;
29819: waveform_sig_loopback =8001;
29820: waveform_sig_loopback =6832;
29821: waveform_sig_loopback =7152;
29822: waveform_sig_loopback =6889;
29823: waveform_sig_loopback =8114;
29824: waveform_sig_loopback =6205;
29825: waveform_sig_loopback =7171;
29826: waveform_sig_loopback =7798;
29827: waveform_sig_loopback =6822;
29828: waveform_sig_loopback =6640;
29829: waveform_sig_loopback =7725;
29830: waveform_sig_loopback =7611;
29831: waveform_sig_loopback =5669;
29832: waveform_sig_loopback =7781;
29833: waveform_sig_loopback =8238;
29834: waveform_sig_loopback =5415;
29835: waveform_sig_loopback =7060;
29836: waveform_sig_loopback =8527;
29837: waveform_sig_loopback =6408;
29838: waveform_sig_loopback =6044;
29839: waveform_sig_loopback =7991;
29840: waveform_sig_loopback =7450;
29841: waveform_sig_loopback =6312;
29842: waveform_sig_loopback =8701;
29843: waveform_sig_loopback =4097;
29844: waveform_sig_loopback =7100;
29845: waveform_sig_loopback =9311;
29846: waveform_sig_loopback =6448;
29847: waveform_sig_loopback =5862;
29848: waveform_sig_loopback =6161;
29849: waveform_sig_loopback =8259;
29850: waveform_sig_loopback =7803;
29851: waveform_sig_loopback =5441;
29852: waveform_sig_loopback =7015;
29853: waveform_sig_loopback =7130;
29854: waveform_sig_loopback =6791;
29855: waveform_sig_loopback =7319;
29856: waveform_sig_loopback =5505;
29857: waveform_sig_loopback =8129;
29858: waveform_sig_loopback =6553;
29859: waveform_sig_loopback =6162;
29860: waveform_sig_loopback =7382;
29861: waveform_sig_loopback =6422;
29862: waveform_sig_loopback =6835;
29863: waveform_sig_loopback =6310;
29864: waveform_sig_loopback =7694;
29865: waveform_sig_loopback =5785;
29866: waveform_sig_loopback =6538;
29867: waveform_sig_loopback =7402;
29868: waveform_sig_loopback =6314;
29869: waveform_sig_loopback =5903;
29870: waveform_sig_loopback =7526;
29871: waveform_sig_loopback =6803;
29872: waveform_sig_loopback =5071;
29873: waveform_sig_loopback =7555;
29874: waveform_sig_loopback =7219;
29875: waveform_sig_loopback =4999;
29876: waveform_sig_loopback =6660;
29877: waveform_sig_loopback =7593;
29878: waveform_sig_loopback =6104;
29879: waveform_sig_loopback =5200;
29880: waveform_sig_loopback =7385;
29881: waveform_sig_loopback =7004;
29882: waveform_sig_loopback =5280;
29883: waveform_sig_loopback =8281;
29884: waveform_sig_loopback =3302;
29885: waveform_sig_loopback =6360;
29886: waveform_sig_loopback =8901;
29887: waveform_sig_loopback =5342;
29888: waveform_sig_loopback =5176;
29889: waveform_sig_loopback =5732;
29890: waveform_sig_loopback =7201;
29891: waveform_sig_loopback =7166;
29892: waveform_sig_loopback =4690;
29893: waveform_sig_loopback =6088;
29894: waveform_sig_loopback =6536;
29895: waveform_sig_loopback =5881;
29896: waveform_sig_loopback =6345;
29897: waveform_sig_loopback =4999;
29898: waveform_sig_loopback =7055;
29899: waveform_sig_loopback =5684;
29900: waveform_sig_loopback =5495;
29901: waveform_sig_loopback =6247;
29902: waveform_sig_loopback =5725;
29903: waveform_sig_loopback =5822;
29904: waveform_sig_loopback =5374;
29905: waveform_sig_loopback =6928;
29906: waveform_sig_loopback =4702;
29907: waveform_sig_loopback =5599;
29908: waveform_sig_loopback =6699;
29909: waveform_sig_loopback =5053;
29910: waveform_sig_loopback =5006;
29911: waveform_sig_loopback =6787;
29912: waveform_sig_loopback =5307;
29913: waveform_sig_loopback =4470;
29914: waveform_sig_loopback =6545;
29915: waveform_sig_loopback =5887;
29916: waveform_sig_loopback =4378;
29917: waveform_sig_loopback =5271;
29918: waveform_sig_loopback =6672;
29919: waveform_sig_loopback =5089;
29920: waveform_sig_loopback =3734;
29921: waveform_sig_loopback =6853;
29922: waveform_sig_loopback =5497;
29923: waveform_sig_loopback =4191;
29924: waveform_sig_loopback =7415;
29925: waveform_sig_loopback =1588;
29926: waveform_sig_loopback =5789;
29927: waveform_sig_loopback =7623;
29928: waveform_sig_loopback =3847;
29929: waveform_sig_loopback =4383;
29930: waveform_sig_loopback =4384;
29931: waveform_sig_loopback =6081;
29932: waveform_sig_loopback =6038;
29933: waveform_sig_loopback =3243;
29934: waveform_sig_loopback =5098;
29935: waveform_sig_loopback =5246;
29936: waveform_sig_loopback =4585;
29937: waveform_sig_loopback =5093;
29938: waveform_sig_loopback =3800;
29939: waveform_sig_loopback =5696;
29940: waveform_sig_loopback =4441;
29941: waveform_sig_loopback =4314;
29942: waveform_sig_loopback =4732;
29943: waveform_sig_loopback =4796;
29944: waveform_sig_loopback =4240;
29945: waveform_sig_loopback =4057;
29946: waveform_sig_loopback =5925;
29947: waveform_sig_loopback =2801;
29948: waveform_sig_loopback =4766;
29949: waveform_sig_loopback =5206;
29950: waveform_sig_loopback =3369;
29951: waveform_sig_loopback =4243;
29952: waveform_sig_loopback =4901;
29953: waveform_sig_loopback =4110;
29954: waveform_sig_loopback =3259;
29955: waveform_sig_loopback =4739;
29956: waveform_sig_loopback =4909;
29957: waveform_sig_loopback =2639;
29958: waveform_sig_loopback =3928;
29959: waveform_sig_loopback =5520;
29960: waveform_sig_loopback =3177;
29961: waveform_sig_loopback =2611;
29962: waveform_sig_loopback =5498;
29963: waveform_sig_loopback =3654;
29964: waveform_sig_loopback =3151;
29965: waveform_sig_loopback =5656;
29966: waveform_sig_loopback =12;
29967: waveform_sig_loopback =4708;
29968: waveform_sig_loopback =5777;
29969: waveform_sig_loopback =2379;
29970: waveform_sig_loopback =2895;
29971: waveform_sig_loopback =2734;
29972: waveform_sig_loopback =4680;
29973: waveform_sig_loopback =4533;
29974: waveform_sig_loopback =1438;
29975: waveform_sig_loopback =3798;
29976: waveform_sig_loopback =3577;
29977: waveform_sig_loopback =2937;
29978: waveform_sig_loopback =3770;
29979: waveform_sig_loopback =1895;
29980: waveform_sig_loopback =4266;
29981: waveform_sig_loopback =2994;
29982: waveform_sig_loopback =2376;
29983: waveform_sig_loopback =3386;
29984: waveform_sig_loopback =3118;
29985: waveform_sig_loopback =2346;
29986: waveform_sig_loopback =2983;
29987: waveform_sig_loopback =3818;
29988: waveform_sig_loopback =1256;
29989: waveform_sig_loopback =3432;
29990: waveform_sig_loopback =3046;
29991: waveform_sig_loopback =2178;
29992: waveform_sig_loopback =2301;
29993: waveform_sig_loopback =3171;
29994: waveform_sig_loopback =2813;
29995: waveform_sig_loopback =1205;
29996: waveform_sig_loopback =3323;
29997: waveform_sig_loopback =3101;
29998: waveform_sig_loopback =762;
29999: waveform_sig_loopback =2626;
30000: waveform_sig_loopback =3608;
30001: waveform_sig_loopback =1341;
30002: waveform_sig_loopback =1046;
30003: waveform_sig_loopback =3711;
30004: waveform_sig_loopback =1844;
30005: waveform_sig_loopback =1811;
30006: waveform_sig_loopback =3498;
30007: waveform_sig_loopback =-1866;
30008: waveform_sig_loopback =3462;
30009: waveform_sig_loopback =3736;
30010: waveform_sig_loopback =770;
30011: waveform_sig_loopback =1034;
30012: waveform_sig_loopback =867;
30013: waveform_sig_loopback =3390;
30014: waveform_sig_loopback =2315;
30015: waveform_sig_loopback =-275;
30016: waveform_sig_loopback =2380;
30017: waveform_sig_loopback =1210;
30018: waveform_sig_loopback =1608;
30019: waveform_sig_loopback =1822;
30020: waveform_sig_loopback =-102;
30021: waveform_sig_loopback =2912;
30022: waveform_sig_loopback =650;
30023: waveform_sig_loopback =762;
30024: waveform_sig_loopback =1822;
30025: waveform_sig_loopback =907;
30026: waveform_sig_loopback =890;
30027: waveform_sig_loopback =999;
30028: waveform_sig_loopback =1817;
30029: waveform_sig_loopback =-110;
30030: waveform_sig_loopback =1236;
30031: waveform_sig_loopback =1344;
30032: waveform_sig_loopback =441;
30033: waveform_sig_loopback =175;
30034: waveform_sig_loopback =1794;
30035: waveform_sig_loopback =615;
30036: waveform_sig_loopback =-651;
30037: waveform_sig_loopback =1640;
30038: waveform_sig_loopback =1058;
30039: waveform_sig_loopback =-913;
30040: waveform_sig_loopback =754;
30041: waveform_sig_loopback =1739;
30042: waveform_sig_loopback =-588;
30043: waveform_sig_loopback =-472;
30044: waveform_sig_loopback =1646;
30045: waveform_sig_loopback =-127;
30046: waveform_sig_loopback =226;
30047: waveform_sig_loopback =1261;
30048: waveform_sig_loopback =-3309;
30049: waveform_sig_loopback =1480;
30050: waveform_sig_loopback =1667;
30051: waveform_sig_loopback =-748;
30052: waveform_sig_loopback =-1250;
30053: waveform_sig_loopback =-570;
30054: waveform_sig_loopback =1501;
30055: waveform_sig_loopback =61;
30056: waveform_sig_loopback =-1689;
30057: waveform_sig_loopback =193;
30058: waveform_sig_loopback =-470;
30059: waveform_sig_loopback =-38;
30060: waveform_sig_loopback =-585;
30061: waveform_sig_loopback =-1456;
30062: waveform_sig_loopback =909;
30063: waveform_sig_loopback =-1363;
30064: waveform_sig_loopback =-782;
30065: waveform_sig_loopback =-467;
30066: waveform_sig_loopback =-722;
30067: waveform_sig_loopback =-1067;
30068: waveform_sig_loopback =-911;
30069: waveform_sig_loopback =43;
30070: waveform_sig_loopback =-2081;
30071: waveform_sig_loopback =-583;
30072: waveform_sig_loopback =-529;
30073: waveform_sig_loopback =-1428;
30074: waveform_sig_loopback =-1721;
30075: waveform_sig_loopback =35;
30076: waveform_sig_loopback =-1445;
30077: waveform_sig_loopback =-2478;
30078: waveform_sig_loopback =144;
30079: waveform_sig_loopback =-1312;
30080: waveform_sig_loopback =-2593;
30081: waveform_sig_loopback =-1038;
30082: waveform_sig_loopback =-515;
30083: waveform_sig_loopback =-2041;
30084: waveform_sig_loopback =-2720;
30085: waveform_sig_loopback =55;
30086: waveform_sig_loopback =-2218;
30087: waveform_sig_loopback =-1787;
30088: waveform_sig_loopback =-283;
30089: waveform_sig_loopback =-5402;
30090: waveform_sig_loopback =-326;
30091: waveform_sig_loopback =-195;
30092: waveform_sig_loopback =-2696;
30093: waveform_sig_loopback =-3062;
30094: waveform_sig_loopback =-2345;
30095: waveform_sig_loopback =-722;
30096: waveform_sig_loopback =-1526;
30097: waveform_sig_loopback =-3573;
30098: waveform_sig_loopback =-1911;
30099: waveform_sig_loopback =-2051;
30100: waveform_sig_loopback =-2094;
30101: waveform_sig_loopback =-2377;
30102: waveform_sig_loopback =-3241;
30103: waveform_sig_loopback =-1222;
30104: waveform_sig_loopback =-2964;
30105: waveform_sig_loopback =-2616;
30106: waveform_sig_loopback =-2463;
30107: waveform_sig_loopback =-2424;
30108: waveform_sig_loopback =-3019;
30109: waveform_sig_loopback =-2727;
30110: waveform_sig_loopback =-1802;
30111: waveform_sig_loopback =-4058;
30112: waveform_sig_loopback =-2285;
30113: waveform_sig_loopback =-2269;
30114: waveform_sig_loopback =-3600;
30115: waveform_sig_loopback =-3299;
30116: waveform_sig_loopback =-1776;
30117: waveform_sig_loopback =-3670;
30118: waveform_sig_loopback =-3884;
30119: waveform_sig_loopback =-1863;
30120: waveform_sig_loopback =-3172;
30121: waveform_sig_loopback =-4197;
30122: waveform_sig_loopback =-3086;
30123: waveform_sig_loopback =-2018;
30124: waveform_sig_loopback =-4069;
30125: waveform_sig_loopback =-4589;
30126: waveform_sig_loopback =-1335;
30127: waveform_sig_loopback =-4251;
30128: waveform_sig_loopback =-3276;
30129: waveform_sig_loopback =-2290;
30130: waveform_sig_loopback =-7403;
30131: waveform_sig_loopback =-1466;
30132: waveform_sig_loopback =-2182;
30133: waveform_sig_loopback =-4757;
30134: waveform_sig_loopback =-4550;
30135: waveform_sig_loopback =-4025;
30136: waveform_sig_loopback =-2323;
30137: waveform_sig_loopback =-3404;
30138: waveform_sig_loopback =-5474;
30139: waveform_sig_loopback =-3294;
30140: waveform_sig_loopback =-3776;
30141: waveform_sig_loopback =-3993;
30142: waveform_sig_loopback =-3958;
30143: waveform_sig_loopback =-4810;
30144: waveform_sig_loopback =-2985;
30145: waveform_sig_loopback =-4622;
30146: waveform_sig_loopback =-4413;
30147: waveform_sig_loopback =-4070;
30148: waveform_sig_loopback =-3932;
30149: waveform_sig_loopback =-5017;
30150: waveform_sig_loopback =-4072;
30151: waveform_sig_loopback =-3452;
30152: waveform_sig_loopback =-5966;
30153: waveform_sig_loopback =-3589;
30154: waveform_sig_loopback =-4144;
30155: waveform_sig_loopback =-5138;
30156: waveform_sig_loopback =-4599;
30157: waveform_sig_loopback =-3758;
30158: waveform_sig_loopback =-5031;
30159: waveform_sig_loopback =-5503;
30160: waveform_sig_loopback =-3606;
30161: waveform_sig_loopback =-4550;
30162: waveform_sig_loopback =-6061;
30163: waveform_sig_loopback =-4392;
30164: waveform_sig_loopback =-3527;
30165: waveform_sig_loopback =-5908;
30166: waveform_sig_loopback =-5836;
30167: waveform_sig_loopback =-2927;
30168: waveform_sig_loopback =-5996;
30169: waveform_sig_loopback =-4573;
30170: waveform_sig_loopback =-3999;
30171: waveform_sig_loopback =-8878;
30172: waveform_sig_loopback =-2714;
30173: waveform_sig_loopback =-3930;
30174: waveform_sig_loopback =-6303;
30175: waveform_sig_loopback =-5876;
30176: waveform_sig_loopback =-5658;
30177: waveform_sig_loopback =-3604;
30178: waveform_sig_loopback =-4874;
30179: waveform_sig_loopback =-7165;
30180: waveform_sig_loopback =-4351;
30181: waveform_sig_loopback =-5527;
30182: waveform_sig_loopback =-5358;
30183: waveform_sig_loopback =-5230;
30184: waveform_sig_loopback =-6536;
30185: waveform_sig_loopback =-4060;
30186: waveform_sig_loopback =-6111;
30187: waveform_sig_loopback =-5912;
30188: waveform_sig_loopback =-5132;
30189: waveform_sig_loopback =-5570;
30190: waveform_sig_loopback =-6289;
30191: waveform_sig_loopback =-5240;
30192: waveform_sig_loopback =-5135;
30193: waveform_sig_loopback =-7017;
30194: waveform_sig_loopback =-4982;
30195: waveform_sig_loopback =-5581;
30196: waveform_sig_loopback =-6368;
30197: waveform_sig_loopback =-6025;
30198: waveform_sig_loopback =-5008;
30199: waveform_sig_loopback =-6299;
30200: waveform_sig_loopback =-6769;
30201: waveform_sig_loopback =-4836;
30202: waveform_sig_loopback =-5736;
30203: waveform_sig_loopback =-7485;
30204: waveform_sig_loopback =-5466;
30205: waveform_sig_loopback =-4767;
30206: waveform_sig_loopback =-7434;
30207: waveform_sig_loopback =-6681;
30208: waveform_sig_loopback =-4283;
30209: waveform_sig_loopback =-7314;
30210: waveform_sig_loopback =-5328;
30211: waveform_sig_loopback =-5762;
30212: waveform_sig_loopback =-9722;
30213: waveform_sig_loopback =-3648;
30214: waveform_sig_loopback =-5484;
30215: waveform_sig_loopback =-7095;
30216: waveform_sig_loopback =-7245;
30217: waveform_sig_loopback =-6747;
30218: waveform_sig_loopback =-4454;
30219: waveform_sig_loopback =-6453;
30220: waveform_sig_loopback =-8005;
30221: waveform_sig_loopback =-5364;
30222: waveform_sig_loopback =-6883;
30223: waveform_sig_loopback =-5999;
30224: waveform_sig_loopback =-6640;
30225: waveform_sig_loopback =-7492;
30226: waveform_sig_loopback =-4882;
30227: waveform_sig_loopback =-7540;
30228: waveform_sig_loopback =-6636;
30229: waveform_sig_loopback =-6202;
30230: waveform_sig_loopback =-6696;
30231: waveform_sig_loopback =-7107;
30232: waveform_sig_loopback =-6215;
30233: waveform_sig_loopback =-6223;
30234: waveform_sig_loopback =-7796;
30235: waveform_sig_loopback =-5962;
30236: waveform_sig_loopback =-6539;
30237: waveform_sig_loopback =-7154;
30238: waveform_sig_loopback =-7013;
30239: waveform_sig_loopback =-5777;
30240: waveform_sig_loopback =-7215;
30241: waveform_sig_loopback =-7755;
30242: waveform_sig_loopback =-5424;
30243: waveform_sig_loopback =-6822;
30244: waveform_sig_loopback =-8321;
30245: waveform_sig_loopback =-5936;
30246: waveform_sig_loopback =-5917;
30247: waveform_sig_loopback =-8132;
30248: waveform_sig_loopback =-7255;
30249: waveform_sig_loopback =-5320;
30250: waveform_sig_loopback =-7900;
30251: waveform_sig_loopback =-6053;
30252: waveform_sig_loopback =-6795;
30253: waveform_sig_loopback =-10081;
30254: waveform_sig_loopback =-4533;
30255: waveform_sig_loopback =-6190;
30256: waveform_sig_loopback =-7687;
30257: waveform_sig_loopback =-8220;
30258: waveform_sig_loopback =-7048;
30259: waveform_sig_loopback =-5226;
30260: waveform_sig_loopback =-7291;
30261: waveform_sig_loopback =-8362;
30262: waveform_sig_loopback =-6236;
30263: waveform_sig_loopback =-7425;
30264: waveform_sig_loopback =-6468;
30265: waveform_sig_loopback =-7555;
30266: waveform_sig_loopback =-7750;
30267: waveform_sig_loopback =-5567;
30268: waveform_sig_loopback =-8201;
30269: waveform_sig_loopback =-6947;
30270: waveform_sig_loopback =-6954;
30271: waveform_sig_loopback =-7161;
30272: waveform_sig_loopback =-7543;
30273: waveform_sig_loopback =-6767;
30274: waveform_sig_loopback =-6773;
30275: waveform_sig_loopback =-8162;
30276: waveform_sig_loopback =-6575;
30277: waveform_sig_loopback =-6869;
30278: waveform_sig_loopback =-7675;
30279: waveform_sig_loopback =-7593;
30280: waveform_sig_loopback =-5902;
30281: waveform_sig_loopback =-8015;
30282: waveform_sig_loopback =-7938;
30283: waveform_sig_loopback =-5702;
30284: waveform_sig_loopback =-7613;
30285: waveform_sig_loopback =-8335;
30286: waveform_sig_loopback =-6426;
30287: waveform_sig_loopback =-6399;
30288: waveform_sig_loopback =-8288;
30289: waveform_sig_loopback =-7763;
30290: waveform_sig_loopback =-5520;
30291: waveform_sig_loopback =-8259;
30292: waveform_sig_loopback =-6352;
30293: waveform_sig_loopback =-7082;
30294: waveform_sig_loopback =-10374;
30295: waveform_sig_loopback =-4718;
30296: waveform_sig_loopback =-6379;
30297: waveform_sig_loopback =-8135;
30298: waveform_sig_loopback =-8364;
30299: waveform_sig_loopback =-7044;
30300: waveform_sig_loopback =-5639;
30301: waveform_sig_loopback =-7445;
30302: waveform_sig_loopback =-8410;
30303: waveform_sig_loopback =-6504;
30304: waveform_sig_loopback =-7426;
30305: waveform_sig_loopback =-6690;
30306: waveform_sig_loopback =-7787;
30307: waveform_sig_loopback =-7495;
30308: waveform_sig_loopback =-6010;
30309: waveform_sig_loopback =-8168;
30310: waveform_sig_loopback =-6871;
30311: waveform_sig_loopback =-7255;
30312: waveform_sig_loopback =-6961;
30313: waveform_sig_loopback =-7769;
30314: waveform_sig_loopback =-6756;
30315: waveform_sig_loopback =-6656;
30316: waveform_sig_loopback =-8415;
30317: waveform_sig_loopback =-6391;
30318: waveform_sig_loopback =-6809;
30319: waveform_sig_loopback =-7861;
30320: waveform_sig_loopback =-7197;
30321: waveform_sig_loopback =-6022;
30322: waveform_sig_loopback =-8085;
30323: waveform_sig_loopback =-7584;
30324: waveform_sig_loopback =-5762;
30325: waveform_sig_loopback =-7587;
30326: waveform_sig_loopback =-8066;
30327: waveform_sig_loopback =-6311;
30328: waveform_sig_loopback =-6276;
30329: waveform_sig_loopback =-8102;
30330: waveform_sig_loopback =-7665;
30331: waveform_sig_loopback =-5172;
30332: waveform_sig_loopback =-8195;
30333: waveform_sig_loopback =-6152;
30334: waveform_sig_loopback =-6805;
30335: waveform_sig_loopback =-10292;
30336: waveform_sig_loopback =-4267;
30337: waveform_sig_loopback =-6113;
30338: waveform_sig_loopback =-8239;
30339: waveform_sig_loopback =-7710;
30340: waveform_sig_loopback =-6849;
30341: waveform_sig_loopback =-5471;
30342: waveform_sig_loopback =-6883;
30343: waveform_sig_loopback =-8400;
30344: waveform_sig_loopback =-5911;
30345: waveform_sig_loopback =-7147;
30346: waveform_sig_loopback =-6508;
30347: waveform_sig_loopback =-7170;
30348: waveform_sig_loopback =-7262;
30349: waveform_sig_loopback =-5630;
30350: waveform_sig_loopback =-7744;
30351: waveform_sig_loopback =-6516;
30352: waveform_sig_loopback =-6823;
30353: waveform_sig_loopback =-6478;
30354: waveform_sig_loopback =-7396;
30355: waveform_sig_loopback =-6205;
30356: waveform_sig_loopback =-6175;
30357: waveform_sig_loopback =-8040;
30358: waveform_sig_loopback =-5699;
30359: waveform_sig_loopback =-6428;
30360: waveform_sig_loopback =-7533;
30361: waveform_sig_loopback =-6267;
30362: waveform_sig_loopback =-5810;
30363: waveform_sig_loopback =-7475;
30364: waveform_sig_loopback =-6782;
30365: waveform_sig_loopback =-5489;
30366: waveform_sig_loopback =-6737;
30367: waveform_sig_loopback =-7621;
30368: waveform_sig_loopback =-5705;
30369: waveform_sig_loopback =-5434;
30370: waveform_sig_loopback =-7836;
30371: waveform_sig_loopback =-6739;
30372: waveform_sig_loopback =-4461;
30373: waveform_sig_loopback =-7825;
30374: waveform_sig_loopback =-5045;
30375: waveform_sig_loopback =-6499;
30376: waveform_sig_loopback =-9541;
30377: waveform_sig_loopback =-3127;
30378: waveform_sig_loopback =-5810;
30379: waveform_sig_loopback =-7399;
30380: waveform_sig_loopback =-6824;
30381: waveform_sig_loopback =-6357;
30382: waveform_sig_loopback =-4355;
30383: waveform_sig_loopback =-6311;
30384: waveform_sig_loopback =-7709;
30385: waveform_sig_loopback =-4818;
30386: waveform_sig_loopback =-6643;
30387: waveform_sig_loopback =-5446;
30388: waveform_sig_loopback =-6400;
30389: waveform_sig_loopback =-6402;
30390: waveform_sig_loopback =-4738;
30391: waveform_sig_loopback =-6873;
30392: waveform_sig_loopback =-5641;
30393: waveform_sig_loopback =-5894;
30394: waveform_sig_loopback =-5504;
30395: waveform_sig_loopback =-6697;
30396: waveform_sig_loopback =-4965;
30397: waveform_sig_loopback =-5446;
30398: waveform_sig_loopback =-7153;
30399: waveform_sig_loopback =-4337;
30400: waveform_sig_loopback =-5896;
30401: waveform_sig_loopback =-6282;
30402: waveform_sig_loopback =-5134;
30403: waveform_sig_loopback =-5152;
30404: waveform_sig_loopback =-6016;
30405: waveform_sig_loopback =-5988;
30406: waveform_sig_loopback =-4356;
30407: waveform_sig_loopback =-5501;
30408: waveform_sig_loopback =-6942;
30409: waveform_sig_loopback =-4141;
30410: waveform_sig_loopback =-4624;
30411: waveform_sig_loopback =-6925;
30412: waveform_sig_loopback =-5165;
30413: waveform_sig_loopback =-3718;
30414: waveform_sig_loopback =-6637;
30415: waveform_sig_loopback =-3688;
30416: waveform_sig_loopback =-5840;
30417: waveform_sig_loopback =-7947;
30418: waveform_sig_loopback =-2038;
30419: waveform_sig_loopback =-4864;
30420: waveform_sig_loopback =-5999;
30421: waveform_sig_loopback =-5823;
30422: waveform_sig_loopback =-5005;
30423: waveform_sig_loopback =-3026;
30424: waveform_sig_loopback =-5399;
30425: waveform_sig_loopback =-6319;
30426: waveform_sig_loopback =-3527;
30427: waveform_sig_loopback =-5477;
30428: waveform_sig_loopback =-4124;
30429: waveform_sig_loopback =-5239;
30430: waveform_sig_loopback =-5183;
30431: waveform_sig_loopback =-3307;
30432: waveform_sig_loopback =-5661;
30433: waveform_sig_loopback =-4716;
30434: waveform_sig_loopback =-4158;
30435: waveform_sig_loopback =-4455;
30436: waveform_sig_loopback =-5328;
30437: waveform_sig_loopback =-3562;
30438: waveform_sig_loopback =-4693;
30439: waveform_sig_loopback =-4993;
30440: waveform_sig_loopback =-3437;
30441: waveform_sig_loopback =-4742;
30442: waveform_sig_loopback =-4487;
30443: waveform_sig_loopback =-4207;
30444: waveform_sig_loopback =-3335;
30445: waveform_sig_loopback =-5021;
30446: waveform_sig_loopback =-4657;
30447: waveform_sig_loopback =-2509;
30448: waveform_sig_loopback =-4664;
30449: waveform_sig_loopback =-5293;
30450: waveform_sig_loopback =-2653;
30451: waveform_sig_loopback =-3367;
30452: waveform_sig_loopback =-5362;
30453: waveform_sig_loopback =-3806;
30454: waveform_sig_loopback =-2274;
30455: waveform_sig_loopback =-5185;
30456: waveform_sig_loopback =-2098;
30457: waveform_sig_loopback =-4754;
30458: waveform_sig_loopback =-6134;
30459: waveform_sig_loopback =-424;
30460: waveform_sig_loopback =-3719;
30461: waveform_sig_loopback =-4243;
30462: waveform_sig_loopback =-4487;
30463: waveform_sig_loopback =-3333;
30464: waveform_sig_loopback =-1427;
30465: waveform_sig_loopback =-4360;
30466: waveform_sig_loopback =-4292;
30467: waveform_sig_loopback =-2161;
30468: waveform_sig_loopback =-4143;
30469: waveform_sig_loopback =-2144;
30470: waveform_sig_loopback =-4116;
30471: waveform_sig_loopback =-3280;
30472: waveform_sig_loopback =-1729;
30473: waveform_sig_loopback =-4487;
30474: waveform_sig_loopback =-2407;
30475: waveform_sig_loopback =-2955;
30476: waveform_sig_loopback =-3043;
30477: waveform_sig_loopback =-3254;
30478: waveform_sig_loopback =-2157;
30479: waveform_sig_loopback =-2888;
30480: waveform_sig_loopback =-3518;
30481: waveform_sig_loopback =-1985;
30482: waveform_sig_loopback =-2602;
30483: waveform_sig_loopback =-3227;
30484: waveform_sig_loopback =-2552;
30485: waveform_sig_loopback =-1527;
30486: waveform_sig_loopback =-3579;
30487: waveform_sig_loopback =-2740;
30488: waveform_sig_loopback =-969;
30489: waveform_sig_loopback =-3115;
30490: waveform_sig_loopback =-3335;
30491: waveform_sig_loopback =-973;
30492: waveform_sig_loopback =-1847;
30493: waveform_sig_loopback =-3555;
30494: waveform_sig_loopback =-1882;
30495: waveform_sig_loopback =-787;
30496: waveform_sig_loopback =-3363;
30497: waveform_sig_loopback =-251;
30498: waveform_sig_loopback =-3321;
30499: waveform_sig_loopback =-3970;
30500: waveform_sig_loopback =979;
30501: waveform_sig_loopback =-1818;
30502: waveform_sig_loopback =-2433;
30503: waveform_sig_loopback =-3104;
30504: waveform_sig_loopback =-972;
30505: waveform_sig_loopback =-41;
30506: waveform_sig_loopback =-2602;
30507: waveform_sig_loopback =-2176;
30508: waveform_sig_loopback =-879;
30509: waveform_sig_loopback =-1817;
30510: waveform_sig_loopback =-610;
30511: waveform_sig_loopback =-2540;
30512: waveform_sig_loopback =-934;
30513: waveform_sig_loopback =-430;
30514: waveform_sig_loopback =-2335;
30515: waveform_sig_loopback =-553;
30516: waveform_sig_loopback =-1420;
30517: waveform_sig_loopback =-775;
30518: waveform_sig_loopback =-1762;
30519: waveform_sig_loopback =-157;
30520: waveform_sig_loopback =-1031;
30521: waveform_sig_loopback =-1827;
30522: waveform_sig_loopback =80;
30523: waveform_sig_loopback =-899;
30524: waveform_sig_loopback =-1337;
30525: waveform_sig_loopback =-615;
30526: waveform_sig_loopback =286;
30527: waveform_sig_loopback =-1791;
30528: waveform_sig_loopback =-745;
30529: waveform_sig_loopback =971;
30530: waveform_sig_loopback =-1566;
30531: waveform_sig_loopback =-1143;
30532: waveform_sig_loopback =766;
30533: waveform_sig_loopback =-155;
30534: waveform_sig_loopback =-1386;
30535: waveform_sig_loopback =-338;
30536: waveform_sig_loopback =1335;
30537: waveform_sig_loopback =-1525;
30538: waveform_sig_loopback =1415;
30539: waveform_sig_loopback =-1254;
30540: waveform_sig_loopback =-2285;
30541: waveform_sig_loopback =3082;
30542: waveform_sig_loopback =130;
30543: waveform_sig_loopback =-1040;
30544: waveform_sig_loopback =-685;
30545: waveform_sig_loopback =767;
30546: waveform_sig_loopback =1677;
30547: waveform_sig_loopback =-399;
30548: waveform_sig_loopback =-632;
30549: waveform_sig_loopback =1230;
30550: waveform_sig_loopback =111;
30551: waveform_sig_loopback =1000;
30552: waveform_sig_loopback =-330;
30553: waveform_sig_loopback =833;
30554: waveform_sig_loopback =1332;
30555: waveform_sig_loopback =-243;
30556: waveform_sig_loopback =1103;
30557: waveform_sig_loopback =632;
30558: waveform_sig_loopback =1035;
30559: waveform_sig_loopback =46;
30560: waveform_sig_loopback =1857;
30561: waveform_sig_loopback =765;
30562: waveform_sig_loopback =41;
30563: waveform_sig_loopback =2039;
30564: waveform_sig_loopback =1029;
30565: waveform_sig_loopback =315;
30566: waveform_sig_loopback =1670;
30567: waveform_sig_loopback =1894;
30568: waveform_sig_loopback =25;
30569: waveform_sig_loopback =1521;
30570: waveform_sig_loopback =2426;
30571: waveform_sig_loopback =642;
30572: waveform_sig_loopback =693;
30573: waveform_sig_loopback =2526;
30574: waveform_sig_loopback =2056;
30575: waveform_sig_loopback =71;
30576: waveform_sig_loopback =1818;
30577: waveform_sig_loopback =3284;
30578: waveform_sig_loopback =-22;
30579: waveform_sig_loopback =3732;
30580: waveform_sig_loopback =240;
30581: waveform_sig_loopback =-297;
30582: waveform_sig_loopback =5287;
30583: waveform_sig_loopback =1526;
30584: waveform_sig_loopback =958;
30585: waveform_sig_loopback =1395;
30586: waveform_sig_loopback =2363;
30587: waveform_sig_loopback =3809;
30588: waveform_sig_loopback =1248;
30589: waveform_sig_loopback =1223;
30590: waveform_sig_loopback =3348;
30591: waveform_sig_loopback =1691;
30592: waveform_sig_loopback =2934;
30593: waveform_sig_loopback =1608;
30594: waveform_sig_loopback =2533;
30595: waveform_sig_loopback =3301;
30596: waveform_sig_loopback =1567;
30597: waveform_sig_loopback =2796;
30598: waveform_sig_loopback =2674;
30599: waveform_sig_loopback =2719;
30600: waveform_sig_loopback =1852;
30601: waveform_sig_loopback =3925;
30602: waveform_sig_loopback =2258;
30603: waveform_sig_loopback =1988;
30604: waveform_sig_loopback =4003;
30605: waveform_sig_loopback =2523;
30606: waveform_sig_loopback =2322;
30607: waveform_sig_loopback =3500;
30608: waveform_sig_loopback =3481;
30609: waveform_sig_loopback =2102;
30610: waveform_sig_loopback =3112;
30611: waveform_sig_loopback =4188;
30612: waveform_sig_loopback =2570;
30613: waveform_sig_loopback =2184;
30614: waveform_sig_loopback =4561;
30615: waveform_sig_loopback =3753;
30616: waveform_sig_loopback =1596;
30617: waveform_sig_loopback =4078;
30618: waveform_sig_loopback =4610;
30619: waveform_sig_loopback =1857;
30620: waveform_sig_loopback =5818;
30621: waveform_sig_loopback =1277;
30622: waveform_sig_loopback =2102;
30623: waveform_sig_loopback =6868;
30624: waveform_sig_loopback =2967;
30625: waveform_sig_loopback =3015;
30626: waveform_sig_loopback =2726;
30627: waveform_sig_loopback =4355;
30628: waveform_sig_loopback =5572;
30629: waveform_sig_loopback =2539;
30630: waveform_sig_loopback =3246;
30631: waveform_sig_loopback =4956;
30632: waveform_sig_loopback =3307;
30633: waveform_sig_loopback =4770;
30634: waveform_sig_loopback =3056;
30635: waveform_sig_loopback =4323;
30636: waveform_sig_loopback =5039;
30637: waveform_sig_loopback =3033;
30638: waveform_sig_loopback =4528;
30639: waveform_sig_loopback =4456;
30640: waveform_sig_loopback =4133;
30641: waveform_sig_loopback =3666;
30642: waveform_sig_loopback =5624;
30643: waveform_sig_loopback =3589;
30644: waveform_sig_loopback =4021;
30645: waveform_sig_loopback =5315;
30646: waveform_sig_loopback =4158;
30647: waveform_sig_loopback =4108;
30648: waveform_sig_loopback =4748;
30649: waveform_sig_loopback =5344;
30650: waveform_sig_loopback =3501;
30651: waveform_sig_loopback =4670;
30652: waveform_sig_loopback =5991;
30653: waveform_sig_loopback =3755;
30654: waveform_sig_loopback =3895;
30655: waveform_sig_loopback =6287;
30656: waveform_sig_loopback =4978;
30657: waveform_sig_loopback =3222;
30658: waveform_sig_loopback =5814;
30659: waveform_sig_loopback =5853;
30660: waveform_sig_loopback =3559;
30661: waveform_sig_loopback =7327;
30662: waveform_sig_loopback =2417;
30663: waveform_sig_loopback =4203;
30664: waveform_sig_loopback =7918;
30665: waveform_sig_loopback =4533;
30666: waveform_sig_loopback =4687;
30667: waveform_sig_loopback =3851;
30668: waveform_sig_loopback =6291;
30669: waveform_sig_loopback =6753;
30670: waveform_sig_loopback =3881;
30671: waveform_sig_loopback =5055;
30672: waveform_sig_loopback =5966;
30673: waveform_sig_loopback =4965;
30674: waveform_sig_loopback =6190;
30675: waveform_sig_loopback =4209;
30676: waveform_sig_loopback =6076;
30677: waveform_sig_loopback =6216;
30678: waveform_sig_loopback =4384;
30679: waveform_sig_loopback =6100;
30680: waveform_sig_loopback =5676;
30681: waveform_sig_loopback =5450;
30682: waveform_sig_loopback =5165;
30683: waveform_sig_loopback =6786;
30684: waveform_sig_loopback =4863;
30685: waveform_sig_loopback =5586;
30686: waveform_sig_loopback =6356;
30687: waveform_sig_loopback =5657;
30688: waveform_sig_loopback =5347;
30689: waveform_sig_loopback =5979;
30690: waveform_sig_loopback =6871;
30691: waveform_sig_loopback =4404;
30692: waveform_sig_loopback =6203;
30693: waveform_sig_loopback =7278;
30694: waveform_sig_loopback =4659;
30695: waveform_sig_loopback =5556;
30696: waveform_sig_loopback =7346;
30697: waveform_sig_loopback =6022;
30698: waveform_sig_loopback =4724;
30699: waveform_sig_loopback =6824;
30700: waveform_sig_loopback =7027;
30701: waveform_sig_loopback =4952;
30702: waveform_sig_loopback =8210;
30703: waveform_sig_loopback =3673;
30704: waveform_sig_loopback =5427;
30705: waveform_sig_loopback =8991;
30706: waveform_sig_loopback =5779;
30707: waveform_sig_loopback =5509;
30708: waveform_sig_loopback =5175;
30709: waveform_sig_loopback =7485;
30710: waveform_sig_loopback =7615;
30711: waveform_sig_loopback =5036;
30712: waveform_sig_loopback =6190;
30713: waveform_sig_loopback =6931;
30714: waveform_sig_loopback =6122;
30715: waveform_sig_loopback =7190;
30716: waveform_sig_loopback =5141;
30717: waveform_sig_loopback =7366;
30718: waveform_sig_loopback =6913;
30719: waveform_sig_loopback =5497;
30720: waveform_sig_loopback =7248;
30721: waveform_sig_loopback =6326;
30722: waveform_sig_loopback =6636;
30723: waveform_sig_loopback =6101;
30724: waveform_sig_loopback =7575;
30725: waveform_sig_loopback =6038;
30726: waveform_sig_loopback =6241;
30727: waveform_sig_loopback =7436;
30728: waveform_sig_loopback =6690;
30729: waveform_sig_loopback =5868;
30730: waveform_sig_loopback =7290;
30731: waveform_sig_loopback =7541;
30732: waveform_sig_loopback =5220;
30733: waveform_sig_loopback =7399;
30734: waveform_sig_loopback =7761;
30735: waveform_sig_loopback =5601;
30736: waveform_sig_loopback =6584;
30737: waveform_sig_loopback =7924;
30738: waveform_sig_loopback =6968;
30739: waveform_sig_loopback =5439;
30740: waveform_sig_loopback =7691;
30741: waveform_sig_loopback =7852;
30742: waveform_sig_loopback =5624;
30743: waveform_sig_loopback =9046;
30744: waveform_sig_loopback =4348;
30745: waveform_sig_loopback =6265;
30746: waveform_sig_loopback =9756;
30747: waveform_sig_loopback =6479;
30748: waveform_sig_loopback =6048;
30749: waveform_sig_loopback =6140;
30750: waveform_sig_loopback =8114;
30751: waveform_sig_loopback =8199;
30752: waveform_sig_loopback =5852;
30753: waveform_sig_loopback =6767;
30754: waveform_sig_loopback =7601;
30755: waveform_sig_loopback =6898;
30756: waveform_sig_loopback =7597;
30757: waveform_sig_loopback =5907;
30758: waveform_sig_loopback =8058;
30759: waveform_sig_loopback =7250;
30760: waveform_sig_loopback =6399;
30761: waveform_sig_loopback =7627;
30762: waveform_sig_loopback =6919;
30763: waveform_sig_loopback =7396;
30764: waveform_sig_loopback =6351;
30765: waveform_sig_loopback =8391;
30766: waveform_sig_loopback =6483;
30767: waveform_sig_loopback =6611;
30768: waveform_sig_loopback =8268;
30769: waveform_sig_loopback =6780;
30770: waveform_sig_loopback =6488;
30771: waveform_sig_loopback =7994;
30772: waveform_sig_loopback =7489;
30773: waveform_sig_loopback =5990;
30774: waveform_sig_loopback =7780;
30775: waveform_sig_loopback =8081;
30776: waveform_sig_loopback =6127;
30777: waveform_sig_loopback =6789;
30778: waveform_sig_loopback =8481;
30779: waveform_sig_loopback =7196;
30780: waveform_sig_loopback =5766;
30781: waveform_sig_loopback =8174;
30782: waveform_sig_loopback =7880;
30783: waveform_sig_loopback =5943;
30784: waveform_sig_loopback =9466;
30785: waveform_sig_loopback =4483;
30786: waveform_sig_loopback =6476;
30787: waveform_sig_loopback =10057;
30788: waveform_sig_loopback =6753;
30789: waveform_sig_loopback =6150;
30790: waveform_sig_loopback =6570;
30791: waveform_sig_loopback =7937;
30792: waveform_sig_loopback =8665;
30793: waveform_sig_loopback =6056;
30794: waveform_sig_loopback =6607;
30795: waveform_sig_loopback =8119;
30796: waveform_sig_loopback =6810;
30797: waveform_sig_loopback =7786;
30798: waveform_sig_loopback =6161;
30799: waveform_sig_loopback =7829;
30800: waveform_sig_loopback =7627;
30801: waveform_sig_loopback =6384;
30802: waveform_sig_loopback =7474;
30803: waveform_sig_loopback =7259;
30804: waveform_sig_loopback =7159;
30805: waveform_sig_loopback =6558;
30806: waveform_sig_loopback =8429;
30807: waveform_sig_loopback =6199;
30808: waveform_sig_loopback =6946;
30809: waveform_sig_loopback =8106;
30810: waveform_sig_loopback =6618;
30811: waveform_sig_loopback =6594;
30812: waveform_sig_loopback =7975;
30813: waveform_sig_loopback =7304;
30814: waveform_sig_loopback =5939;
30815: waveform_sig_loopback =7746;
30816: waveform_sig_loopback =7845;
30817: waveform_sig_loopback =6124;
30818: waveform_sig_loopback =6556;
30819: waveform_sig_loopback =8448;
30820: waveform_sig_loopback =7054;
30821: waveform_sig_loopback =5318;
30822: waveform_sig_loopback =8375;
30823: waveform_sig_loopback =7551;
30824: waveform_sig_loopback =5756;
30825: waveform_sig_loopback =9383;
30826: waveform_sig_loopback =3737;
30827: waveform_sig_loopback =6905;
30828: waveform_sig_loopback =9795;
30829: waveform_sig_loopback =5905;
30830: waveform_sig_loopback =6261;
30831: waveform_sig_loopback =6181;
30832: waveform_sig_loopback =7816;
30833: waveform_sig_loopback =8381;
30834: waveform_sig_loopback =5263;
30835: waveform_sig_loopback =6821;
30836: waveform_sig_loopback =7622;
30837: waveform_sig_loopback =6249;
30838: waveform_sig_loopback =7631;
30839: waveform_sig_loopback =5598;
30840: waveform_sig_loopback =7618;
30841: waveform_sig_loopback =7134;
30842: waveform_sig_loopback =5860;
30843: waveform_sig_loopback =7284;
30844: waveform_sig_loopback =6795;
30845: waveform_sig_loopback =6552;
30846: waveform_sig_loopback =6253;
30847: waveform_sig_loopback =7969;
30848: waveform_sig_loopback =5554;
30849: waveform_sig_loopback =6607;
30850: waveform_sig_loopback =7558;
30851: waveform_sig_loopback =5998;
30852: waveform_sig_loopback =6293;
30853: waveform_sig_loopback =7202;
30854: waveform_sig_loopback =6735;
30855: waveform_sig_loopback =5587;
30856: waveform_sig_loopback =6906;
30857: waveform_sig_loopback =7537;
30858: waveform_sig_loopback =5304;
30859: waveform_sig_loopback =5969;
30860: waveform_sig_loopback =8174;
30861: waveform_sig_loopback =5910;
30862: waveform_sig_loopback =5004;
30863: waveform_sig_loopback =7858;
30864: waveform_sig_loopback =6454;
30865: waveform_sig_loopback =5596;
30866: waveform_sig_loopback =8393;
30867: waveform_sig_loopback =2907;
30868: waveform_sig_loopback =6710;
30869: waveform_sig_loopback =8617;
30870: waveform_sig_loopback =5436;
30871: waveform_sig_loopback =5504;
30872: waveform_sig_loopback =5183;
30873: waveform_sig_loopback =7474;
30874: waveform_sig_loopback =7313;
30875: waveform_sig_loopback =4397;
30876: waveform_sig_loopback =6274;
30877: waveform_sig_loopback =6487;
30878: waveform_sig_loopback =5682;
30879: waveform_sig_loopback =6745;
30880: waveform_sig_loopback =4591;
30881: waveform_sig_loopback =7029;
30882: waveform_sig_loopback =6096;
30883: waveform_sig_loopback =5055;
30884: waveform_sig_loopback =6407;
30885: waveform_sig_loopback =5914;
30886: waveform_sig_loopback =5528;
30887: waveform_sig_loopback =5560;
30888: waveform_sig_loopback =6923;
30889: waveform_sig_loopback =4508;
30890: waveform_sig_loopback =6084;
30891: waveform_sig_loopback =6158;
30892: waveform_sig_loopback =5317;
30893: waveform_sig_loopback =5277;
30894: waveform_sig_loopback =6022;
30895: waveform_sig_loopback =6153;
30896: waveform_sig_loopback =4118;
30897: waveform_sig_loopback =6220;
30898: waveform_sig_loopback =6536;
30899: waveform_sig_loopback =3840;
30900: waveform_sig_loopback =5462;
30901: waveform_sig_loopback =6797;
30902: waveform_sig_loopback =4808;
30903: waveform_sig_loopback =4191;
30904: waveform_sig_loopback =6484;
30905: waveform_sig_loopback =5513;
30906: waveform_sig_loopback =4529;
30907: waveform_sig_loopback =7111;
30908: waveform_sig_loopback =1838;
30909: waveform_sig_loopback =5680;
30910: waveform_sig_loopback =7481;
30911: waveform_sig_loopback =4164;
30912: waveform_sig_loopback =4301;
30913: waveform_sig_loopback =4096;
30914: waveform_sig_loopback =6310;
30915: waveform_sig_loopback =6067;
30916: waveform_sig_loopback =3043;
30917: waveform_sig_loopback =5352;
30918: waveform_sig_loopback =4984;
30919: waveform_sig_loopback =4603;
30920: waveform_sig_loopback =5531;
30921: waveform_sig_loopback =3106;
30922: waveform_sig_loopback =6175;
30923: waveform_sig_loopback =4471;
30924: waveform_sig_loopback =3817;
30925: waveform_sig_loopback =5407;
30926: waveform_sig_loopback =4190;
30927: waveform_sig_loopback =4534;
30928: waveform_sig_loopback =4228;
30929: waveform_sig_loopback =5310;
30930: waveform_sig_loopback =3582;
30931: waveform_sig_loopback =4325;
30932: waveform_sig_loopback =5028;
30933: waveform_sig_loopback =3944;
30934: waveform_sig_loopback =3674;
30935: waveform_sig_loopback =5114;
30936: waveform_sig_loopback =4315;
30937: waveform_sig_loopback =2833;
30938: waveform_sig_loopback =4977;
30939: waveform_sig_loopback =4914;
30940: waveform_sig_loopback =2519;
30941: waveform_sig_loopback =4081;
30942: waveform_sig_loopback =5338;
30943: waveform_sig_loopback =3263;
30944: waveform_sig_loopback =2912;
30945: waveform_sig_loopback =4998;
30946: waveform_sig_loopback =3961;
30947: waveform_sig_loopback =3189;
30948: waveform_sig_loopback =5418;
30949: waveform_sig_loopback =468;
30950: waveform_sig_loopback =4268;
30951: waveform_sig_loopback =5821;
30952: waveform_sig_loopback =2843;
30953: waveform_sig_loopback =2538;
30954: waveform_sig_loopback =2806;
30955: waveform_sig_loopback =4925;
30956: waveform_sig_loopback =4147;
30957: waveform_sig_loopback =1863;
30958: waveform_sig_loopback =3705;
30959: waveform_sig_loopback =3339;
30960: waveform_sig_loopback =3409;
30961: waveform_sig_loopback =3459;
30962: waveform_sig_loopback =1935;
30963: waveform_sig_loopback =4613;
30964: waveform_sig_loopback =2486;
30965: waveform_sig_loopback =2809;
30966: waveform_sig_loopback =3355;
30967: waveform_sig_loopback =2753;
30968: waveform_sig_loopback =3014;
30969: waveform_sig_loopback =2353;
30970: waveform_sig_loopback =4010;
30971: waveform_sig_loopback =1681;
30972: waveform_sig_loopback =2734;
30973: waveform_sig_loopback =3558;
30974: waveform_sig_loopback =2035;
30975: waveform_sig_loopback =2135;
30976: waveform_sig_loopback =3486;
30977: waveform_sig_loopback =2514;
30978: waveform_sig_loopback =1264;
30979: waveform_sig_loopback =3425;
30980: waveform_sig_loopback =2990;
30981: waveform_sig_loopback =890;
30982: waveform_sig_loopback =2551;
30983: waveform_sig_loopback =3407;
30984: waveform_sig_loopback =1604;
30985: waveform_sig_loopback =1111;
30986: waveform_sig_loopback =3262;
30987: waveform_sig_loopback =2320;
30988: waveform_sig_loopback =1325;
30989: waveform_sig_loopback =3644;
30990: waveform_sig_loopback =-1212;
30991: waveform_sig_loopback =2504;
30992: waveform_sig_loopback =4269;
30993: waveform_sig_loopback =869;
30994: waveform_sig_loopback =636;
30995: waveform_sig_loopback =1477;
30996: waveform_sig_loopback =2777;
30997: waveform_sig_loopback =2503;
30998: waveform_sig_loopback =121;
30999: waveform_sig_loopback =1672;
31000: waveform_sig_loopback =1905;
31001: waveform_sig_loopback =1358;
31002: waveform_sig_loopback =1618;
31003: waveform_sig_loopback =420;
31004: waveform_sig_loopback =2464;
31005: waveform_sig_loopback =918;
31006: waveform_sig_loopback =936;
31007: waveform_sig_loopback =1391;
31008: waveform_sig_loopback =1203;
31009: waveform_sig_loopback =891;
31010: waveform_sig_loopback =700;
31011: waveform_sig_loopback =2178;
31012: waveform_sig_loopback =-281;
31013: waveform_sig_loopback =1073;
31014: waveform_sig_loopback =1647;
31015: waveform_sig_loopback =207;
31016: waveform_sig_loopback =276;
31017: waveform_sig_loopback =1839;
31018: waveform_sig_loopback =322;
31019: waveform_sig_loopback =-353;
31020: waveform_sig_loopback =1624;
31021: waveform_sig_loopback =768;
31022: waveform_sig_loopback =-597;
31023: waveform_sig_loopback =470;
31024: waveform_sig_loopback =1623;
31025: waveform_sig_loopback =-112;
31026: waveform_sig_loopback =-1142;
31027: waveform_sig_loopback =1989;
31028: waveform_sig_loopback =31;
31029: waveform_sig_loopback =-462;
31030: waveform_sig_loopback =2067;
31031: waveform_sig_loopback =-3729;
31032: waveform_sig_loopback =1273;
31033: waveform_sig_loopback =2154;
31034: waveform_sig_loopback =-1341;
31035: waveform_sig_loopback =-807;
31036: waveform_sig_loopback =-607;
31037: waveform_sig_loopback =985;
31038: waveform_sig_loopback =681;
31039: waveform_sig_loopback =-2060;
31040: waveform_sig_loopback =99;
31041: waveform_sig_loopback =-43;
31042: waveform_sig_loopback =-696;
31043: waveform_sig_loopback =-134;
31044: waveform_sig_loopback =-1465;
31045: waveform_sig_loopback =435;
31046: waveform_sig_loopback =-855;
31047: waveform_sig_loopback =-1071;
31048: waveform_sig_loopback =-470;
31049: waveform_sig_loopback =-526;
31050: waveform_sig_loopback =-1320;
31051: waveform_sig_loopback =-917;
31052: waveform_sig_loopback =242;
31053: waveform_sig_loopback =-2409;
31054: waveform_sig_loopback =-534;
31055: waveform_sig_loopback =-435;
31056: waveform_sig_loopback =-1816;
31057: waveform_sig_loopback =-1287;
31058: waveform_sig_loopback =-311;
31059: waveform_sig_loopback =-1563;
31060: waveform_sig_loopback =-2043;
31061: waveform_sig_loopback =-479;
31062: waveform_sig_loopback =-907;
31063: waveform_sig_loopback =-2633;
31064: waveform_sig_loopback =-1465;
31065: waveform_sig_loopback =20;
31066: waveform_sig_loopback =-2411;
31067: waveform_sig_loopback =-2815;
31068: waveform_sig_loopback =320;
31069: waveform_sig_loopback =-2318;
31070: waveform_sig_loopback =-1870;
31071: waveform_sig_loopback =-95;
31072: waveform_sig_loopback =-5763;
31073: waveform_sig_loopback =-49;
31074: waveform_sig_loopback =-207;
31075: waveform_sig_loopback =-3131;
31076: waveform_sig_loopback =-2537;
31077: waveform_sig_loopback =-2763;
31078: waveform_sig_loopback =-508;
31079: waveform_sig_loopback =-1425;
31080: waveform_sig_loopback =-4068;
31081: waveform_sig_loopback =-1344;
31082: waveform_sig_loopback =-2235;
31083: waveform_sig_loopback =-2383;
31084: waveform_sig_loopback =-1975;
31085: waveform_sig_loopback =-3537;
31086: waveform_sig_loopback =-1051;
31087: waveform_sig_loopback =-2888;
31088: waveform_sig_loopback =-2912;
31089: waveform_sig_loopback =-2233;
31090: waveform_sig_loopback =-2344;
31091: waveform_sig_loopback =-3259;
31092: waveform_sig_loopback =-2538;
31093: waveform_sig_loopback =-1746;
31094: waveform_sig_loopback =-4269;
31095: waveform_sig_loopback =-1982;
31096: waveform_sig_loopback =-2648;
31097: waveform_sig_loopback =-3334;
31098: waveform_sig_loopback =-3082;
31099: waveform_sig_loopback =-2372;
31100: waveform_sig_loopback =-3052;
31101: waveform_sig_loopback =-4113;
31102: waveform_sig_loopback =-2100;
31103: waveform_sig_loopback =-2610;
31104: waveform_sig_loopback =-4770;
31105: waveform_sig_loopback =-2848;
31106: waveform_sig_loopback =-1852;
31107: waveform_sig_loopback =-4453;
31108: waveform_sig_loopback =-4191;
31109: waveform_sig_loopback =-1666;
31110: waveform_sig_loopback =-4144;
31111: waveform_sig_loopback =-3239;
31112: waveform_sig_loopback =-2345;
31113: waveform_sig_loopback =-7266;
31114: waveform_sig_loopback =-1589;
31115: waveform_sig_loopback =-2265;
31116: waveform_sig_loopback =-4527;
31117: waveform_sig_loopback =-4487;
31118: waveform_sig_loopback =-4511;
31119: waveform_sig_loopback =-1949;
31120: waveform_sig_loopback =-3469;
31121: waveform_sig_loopback =-5595;
31122: waveform_sig_loopback =-2995;
31123: waveform_sig_loopback =-4248;
31124: waveform_sig_loopback =-3656;
31125: waveform_sig_loopback =-3870;
31126: waveform_sig_loopback =-5170;
31127: waveform_sig_loopback =-2464;
31128: waveform_sig_loopback =-4877;
31129: waveform_sig_loopback =-4427;
31130: waveform_sig_loopback =-3746;
31131: waveform_sig_loopback =-4206;
31132: waveform_sig_loopback =-4738;
31133: waveform_sig_loopback =-4312;
31134: waveform_sig_loopback =-3603;
31135: waveform_sig_loopback =-5498;
31136: waveform_sig_loopback =-3742;
31137: waveform_sig_loopback =-4476;
31138: waveform_sig_loopback =-4863;
31139: waveform_sig_loopback =-4800;
31140: waveform_sig_loopback =-3671;
31141: waveform_sig_loopback =-4782;
31142: waveform_sig_loopback =-6115;
31143: waveform_sig_loopback =-3127;
31144: waveform_sig_loopback =-4480;
31145: waveform_sig_loopback =-6461;
31146: waveform_sig_loopback =-4042;
31147: waveform_sig_loopback =-3844;
31148: waveform_sig_loopback =-5743;
31149: waveform_sig_loopback =-5813;
31150: waveform_sig_loopback =-3404;
31151: waveform_sig_loopback =-5465;
31152: waveform_sig_loopback =-4896;
31153: waveform_sig_loopback =-4097;
31154: waveform_sig_loopback =-8537;
31155: waveform_sig_loopback =-3141;
31156: waveform_sig_loopback =-3765;
31157: waveform_sig_loopback =-6061;
31158: waveform_sig_loopback =-6223;
31159: waveform_sig_loopback =-5467;
31160: waveform_sig_loopback =-3580;
31161: waveform_sig_loopback =-5135;
31162: waveform_sig_loopback =-6797;
31163: waveform_sig_loopback =-4571;
31164: waveform_sig_loopback =-5573;
31165: waveform_sig_loopback =-5066;
31166: waveform_sig_loopback =-5522;
31167: waveform_sig_loopback =-6397;
31168: waveform_sig_loopback =-3968;
31169: waveform_sig_loopback =-6388;
31170: waveform_sig_loopback =-5586;
31171: waveform_sig_loopback =-5226;
31172: waveform_sig_loopback =-5725;
31173: waveform_sig_loopback =-5972;
31174: waveform_sig_loopback =-5519;
31175: waveform_sig_loopback =-5033;
31176: waveform_sig_loopback =-6814;
31177: waveform_sig_loopback =-5450;
31178: waveform_sig_loopback =-5305;
31179: waveform_sig_loopback =-6305;
31180: waveform_sig_loopback =-6468;
31181: waveform_sig_loopback =-4540;
31182: waveform_sig_loopback =-6563;
31183: waveform_sig_loopback =-6910;
31184: waveform_sig_loopback =-4517;
31185: waveform_sig_loopback =-6181;
31186: waveform_sig_loopback =-7095;
31187: waveform_sig_loopback =-5602;
31188: waveform_sig_loopback =-5019;
31189: waveform_sig_loopback =-6897;
31190: waveform_sig_loopback =-7139;
31191: waveform_sig_loopback =-4251;
31192: waveform_sig_loopback =-7019;
31193: waveform_sig_loopback =-5867;
31194: waveform_sig_loopback =-5290;
31195: waveform_sig_loopback =-9822;
31196: waveform_sig_loopback =-4045;
31197: waveform_sig_loopback =-5047;
31198: waveform_sig_loopback =-7210;
31199: waveform_sig_loopback =-7363;
31200: waveform_sig_loopback =-6503;
31201: waveform_sig_loopback =-4765;
31202: waveform_sig_loopback =-6301;
31203: waveform_sig_loopback =-7754;
31204: waveform_sig_loopback =-5828;
31205: waveform_sig_loopback =-6462;
31206: waveform_sig_loopback =-6147;
31207: waveform_sig_loopback =-6774;
31208: waveform_sig_loopback =-7070;
31209: waveform_sig_loopback =-5307;
31210: waveform_sig_loopback =-7353;
31211: waveform_sig_loopback =-6485;
31212: waveform_sig_loopback =-6554;
31213: waveform_sig_loopback =-6398;
31214: waveform_sig_loopback =-7137;
31215: waveform_sig_loopback =-6563;
31216: waveform_sig_loopback =-5755;
31217: waveform_sig_loopback =-8126;
31218: waveform_sig_loopback =-6030;
31219: waveform_sig_loopback =-6184;
31220: waveform_sig_loopback =-7536;
31221: waveform_sig_loopback =-6848;
31222: waveform_sig_loopback =-5704;
31223: waveform_sig_loopback =-7516;
31224: waveform_sig_loopback =-7433;
31225: waveform_sig_loopback =-5692;
31226: waveform_sig_loopback =-6859;
31227: waveform_sig_loopback =-8008;
31228: waveform_sig_loopback =-6436;
31229: waveform_sig_loopback =-5685;
31230: waveform_sig_loopback =-7988;
31231: waveform_sig_loopback =-7769;
31232: waveform_sig_loopback =-4955;
31233: waveform_sig_loopback =-7954;
31234: waveform_sig_loopback =-6388;
31235: waveform_sig_loopback =-6267;
31236: waveform_sig_loopback =-10499;
31237: waveform_sig_loopback =-4622;
31238: waveform_sig_loopback =-5850;
31239: waveform_sig_loopback =-8059;
31240: waveform_sig_loopback =-7971;
31241: waveform_sig_loopback =-7058;
31242: waveform_sig_loopback =-5618;
31243: waveform_sig_loopback =-6780;
31244: waveform_sig_loopback =-8591;
31245: waveform_sig_loopback =-6436;
31246: waveform_sig_loopback =-6923;
31247: waveform_sig_loopback =-7054;
31248: waveform_sig_loopback =-7143;
31249: waveform_sig_loopback =-7733;
31250: waveform_sig_loopback =-6064;
31251: waveform_sig_loopback =-7589;
31252: waveform_sig_loopback =-7354;
31253: waveform_sig_loopback =-6996;
31254: waveform_sig_loopback =-6784;
31255: waveform_sig_loopback =-8023;
31256: waveform_sig_loopback =-6549;
31257: waveform_sig_loopback =-6599;
31258: waveform_sig_loopback =-8587;
31259: waveform_sig_loopback =-6144;
31260: waveform_sig_loopback =-7068;
31261: waveform_sig_loopback =-7741;
31262: waveform_sig_loopback =-7300;
31263: waveform_sig_loopback =-6234;
31264: waveform_sig_loopback =-7736;
31265: waveform_sig_loopback =-7946;
31266: waveform_sig_loopback =-5967;
31267: waveform_sig_loopback =-7256;
31268: waveform_sig_loopback =-8372;
31269: waveform_sig_loopback =-6698;
31270: waveform_sig_loopback =-6054;
31271: waveform_sig_loopback =-8362;
31272: waveform_sig_loopback =-7998;
31273: waveform_sig_loopback =-5118;
31274: waveform_sig_loopback =-8555;
31275: waveform_sig_loopback =-6367;
31276: waveform_sig_loopback =-6703;
31277: waveform_sig_loopback =-10926;
31278: waveform_sig_loopback =-4386;
31279: waveform_sig_loopback =-6433;
31280: waveform_sig_loopback =-8372;
31281: waveform_sig_loopback =-7810;
31282: waveform_sig_loopback =-7663;
31283: waveform_sig_loopback =-5448;
31284: waveform_sig_loopback =-7084;
31285: waveform_sig_loopback =-9014;
31286: waveform_sig_loopback =-6011;
31287: waveform_sig_loopback =-7634;
31288: waveform_sig_loopback =-6926;
31289: waveform_sig_loopback =-7193;
31290: waveform_sig_loopback =-8147;
31291: waveform_sig_loopback =-5695;
31292: waveform_sig_loopback =-8036;
31293: waveform_sig_loopback =-7326;
31294: waveform_sig_loopback =-6808;
31295: waveform_sig_loopback =-7114;
31296: waveform_sig_loopback =-7828;
31297: waveform_sig_loopback =-6579;
31298: waveform_sig_loopback =-6759;
31299: waveform_sig_loopback =-8454;
31300: waveform_sig_loopback =-6198;
31301: waveform_sig_loopback =-7057;
31302: waveform_sig_loopback =-7748;
31303: waveform_sig_loopback =-7088;
31304: waveform_sig_loopback =-6366;
31305: waveform_sig_loopback =-7614;
31306: waveform_sig_loopback =-7830;
31307: waveform_sig_loopback =-5994;
31308: waveform_sig_loopback =-6939;
31309: waveform_sig_loopback =-8609;
31310: waveform_sig_loopback =-6239;
31311: waveform_sig_loopback =-5940;
31312: waveform_sig_loopback =-8554;
31313: waveform_sig_loopback =-7316;
31314: waveform_sig_loopback =-5288;
31315: waveform_sig_loopback =-8349;
31316: waveform_sig_loopback =-5809;
31317: waveform_sig_loopback =-7049;
31318: waveform_sig_loopback =-10273;
31319: waveform_sig_loopback =-4121;
31320: waveform_sig_loopback =-6512;
31321: waveform_sig_loopback =-7721;
31322: waveform_sig_loopback =-7936;
31323: waveform_sig_loopback =-7180;
31324: waveform_sig_loopback =-4931;
31325: waveform_sig_loopback =-7234;
31326: waveform_sig_loopback =-8364;
31327: waveform_sig_loopback =-5717;
31328: waveform_sig_loopback =-7432;
31329: waveform_sig_loopback =-6214;
31330: waveform_sig_loopback =-7236;
31331: waveform_sig_loopback =-7539;
31332: waveform_sig_loopback =-5177;
31333: waveform_sig_loopback =-7913;
31334: waveform_sig_loopback =-6684;
31335: waveform_sig_loopback =-6512;
31336: waveform_sig_loopback =-6703;
31337: waveform_sig_loopback =-7326;
31338: waveform_sig_loopback =-6104;
31339: waveform_sig_loopback =-6440;
31340: waveform_sig_loopback =-7772;
31341: waveform_sig_loopback =-5750;
31342: waveform_sig_loopback =-6693;
31343: waveform_sig_loopback =-7009;
31344: waveform_sig_loopback =-6790;
31345: waveform_sig_loopback =-5675;
31346: waveform_sig_loopback =-7068;
31347: waveform_sig_loopback =-7472;
31348: waveform_sig_loopback =-5018;
31349: waveform_sig_loopback =-6729;
31350: waveform_sig_loopback =-8004;
31351: waveform_sig_loopback =-5268;
31352: waveform_sig_loopback =-5773;
31353: waveform_sig_loopback =-7691;
31354: waveform_sig_loopback =-6585;
31355: waveform_sig_loopback =-4917;
31356: waveform_sig_loopback =-7367;
31357: waveform_sig_loopback =-5277;
31358: waveform_sig_loopback =-6584;
31359: waveform_sig_loopback =-9205;
31360: waveform_sig_loopback =-3616;
31361: waveform_sig_loopback =-5647;
31362: waveform_sig_loopback =-7047;
31363: waveform_sig_loopback =-7363;
31364: waveform_sig_loopback =-6093;
31365: waveform_sig_loopback =-4341;
31366: waveform_sig_loopback =-6554;
31367: waveform_sig_loopback =-7404;
31368: waveform_sig_loopback =-5084;
31369: waveform_sig_loopback =-6586;
31370: waveform_sig_loopback =-5250;
31371: waveform_sig_loopback =-6633;
31372: waveform_sig_loopback =-6468;
31373: waveform_sig_loopback =-4427;
31374: waveform_sig_loopback =-7200;
31375: waveform_sig_loopback =-5548;
31376: waveform_sig_loopback =-5722;
31377: waveform_sig_loopback =-5915;
31378: waveform_sig_loopback =-6169;
31379: waveform_sig_loopback =-5314;
31380: waveform_sig_loopback =-5547;
31381: waveform_sig_loopback =-6640;
31382: waveform_sig_loopback =-5109;
31383: waveform_sig_loopback =-5343;
31384: waveform_sig_loopback =-6294;
31385: waveform_sig_loopback =-5789;
31386: waveform_sig_loopback =-4348;
31387: waveform_sig_loopback =-6589;
31388: waveform_sig_loopback =-6013;
31389: waveform_sig_loopback =-4084;
31390: waveform_sig_loopback =-5915;
31391: waveform_sig_loopback =-6617;
31392: waveform_sig_loopback =-4410;
31393: waveform_sig_loopback =-4626;
31394: waveform_sig_loopback =-6618;
31395: waveform_sig_loopback =-5536;
31396: waveform_sig_loopback =-3770;
31397: waveform_sig_loopback =-6340;
31398: waveform_sig_loopback =-4046;
31399: waveform_sig_loopback =-5635;
31400: waveform_sig_loopback =-7927;
31401: waveform_sig_loopback =-2482;
31402: waveform_sig_loopback =-4478;
31403: waveform_sig_loopback =-5964;
31404: waveform_sig_loopback =-6206;
31405: waveform_sig_loopback =-4611;
31406: waveform_sig_loopback =-3383;
31407: waveform_sig_loopback =-5358;
31408: waveform_sig_loopback =-6033;
31409: waveform_sig_loopback =-4082;
31410: waveform_sig_loopback =-5140;
31411: waveform_sig_loopback =-4169;
31412: waveform_sig_loopback =-5536;
31413: waveform_sig_loopback =-4839;
31414: waveform_sig_loopback =-3552;
31415: waveform_sig_loopback =-5762;
31416: waveform_sig_loopback =-4168;
31417: waveform_sig_loopback =-4714;
31418: waveform_sig_loopback =-4305;
31419: waveform_sig_loopback =-5113;
31420: waveform_sig_loopback =-3936;
31421: waveform_sig_loopback =-4080;
31422: waveform_sig_loopback =-5530;
31423: waveform_sig_loopback =-3504;
31424: waveform_sig_loopback =-4075;
31425: waveform_sig_loopback =-5061;
31426: waveform_sig_loopback =-4087;
31427: waveform_sig_loopback =-3122;
31428: waveform_sig_loopback =-5275;
31429: waveform_sig_loopback =-4425;
31430: waveform_sig_loopback =-2788;
31431: waveform_sig_loopback =-4510;
31432: waveform_sig_loopback =-5044;
31433: waveform_sig_loopback =-3046;
31434: waveform_sig_loopback =-3218;
31435: waveform_sig_loopback =-5120;
31436: waveform_sig_loopback =-4103;
31437: waveform_sig_loopback =-2143;
31438: waveform_sig_loopback =-4985;
31439: waveform_sig_loopback =-2547;
31440: waveform_sig_loopback =-4090;
31441: waveform_sig_loopback =-6506;
31442: waveform_sig_loopback =-749;
31443: waveform_sig_loopback =-2995;
31444: waveform_sig_loopback =-4775;
31445: waveform_sig_loopback =-4289;
31446: waveform_sig_loopback =-3200;
31447: waveform_sig_loopback =-1892;
31448: waveform_sig_loopback =-3602;
31449: waveform_sig_loopback =-4723;
31450: waveform_sig_loopback =-2293;
31451: waveform_sig_loopback =-3563;
31452: waveform_sig_loopback =-2766;
31453: waveform_sig_loopback =-3729;
31454: waveform_sig_loopback =-3276;
31455: waveform_sig_loopback =-2040;
31456: waveform_sig_loopback =-3955;
31457: waveform_sig_loopback =-2712;
31458: waveform_sig_loopback =-2978;
31459: waveform_sig_loopback =-2605;
31460: waveform_sig_loopback =-3675;
31461: waveform_sig_loopback =-1996;
31462: waveform_sig_loopback =-2648;
31463: waveform_sig_loopback =-3930;
31464: waveform_sig_loopback =-1633;
31465: waveform_sig_loopback =-2601;
31466: waveform_sig_loopback =-3426;
31467: waveform_sig_loopback =-2253;
31468: waveform_sig_loopback =-1701;
31469: waveform_sig_loopback =-3502;
31470: waveform_sig_loopback =-2589;
31471: waveform_sig_loopback =-1300;
31472: waveform_sig_loopback =-2754;
31473: waveform_sig_loopback =-3379;
31474: waveform_sig_loopback =-1333;
31475: waveform_sig_loopback =-1392;
31476: waveform_sig_loopback =-3664;
31477: waveform_sig_loopback =-2222;
31478: waveform_sig_loopback =-293;
31479: waveform_sig_loopback =-3697;
31480: waveform_sig_loopback =-338;
31481: waveform_sig_loopback =-2773;
31482: waveform_sig_loopback =-4697;
31483: waveform_sig_loopback =1235;
31484: waveform_sig_loopback =-1802;
31485: waveform_sig_loopback =-2694;
31486: waveform_sig_loopback =-2431;
31487: waveform_sig_loopback =-1820;
31488: waveform_sig_loopback =73;
31489: waveform_sig_loopback =-1942;
31490: waveform_sig_loopback =-2919;
31491: waveform_sig_loopback =-381;
31492: waveform_sig_loopback =-2149;
31493: waveform_sig_loopback =-575;
31494: waveform_sig_loopback =-1946;
31495: waveform_sig_loopback =-1717;
31496: waveform_sig_loopback =-82;
31497: waveform_sig_loopback =-2138;
31498: waveform_sig_loopback =-903;
31499: waveform_sig_loopback =-1327;
31500: waveform_sig_loopback =-790;
31501: waveform_sig_loopback =-1765;
31502: waveform_sig_loopback =-81;
31503: waveform_sig_loopback =-1117;
31504: waveform_sig_loopback =-2031;
31505: waveform_sig_loopback =547;
31506: waveform_sig_loopback =-1215;
31507: waveform_sig_loopback =-1398;
31508: waveform_sig_loopback =-289;
31509: waveform_sig_loopback =-166;
31510: waveform_sig_loopback =-1428;
31511: waveform_sig_loopback =-922;
31512: waveform_sig_loopback =703;
31513: waveform_sig_loopback =-979;
31514: waveform_sig_loopback =-1709;
31515: waveform_sig_loopback =895;
31516: waveform_sig_loopback =258;
31517: waveform_sig_loopback =-1975;
31518: waveform_sig_loopback =-23;
31519: waveform_sig_loopback =1378;
31520: waveform_sig_loopback =-1814;
31521: waveform_sig_loopback =1760;
31522: waveform_sig_loopback =-1336;
31523: waveform_sig_loopback =-2507;
31524: waveform_sig_loopback =3296;
31525: waveform_sig_loopback =-150;
31526: waveform_sig_loopback =-709;
31527: waveform_sig_loopback =-745;
31528: waveform_sig_loopback =325;
31529: waveform_sig_loopback =2257;
31530: waveform_sig_loopback =-624;
31531: waveform_sig_loopback =-818;
31532: waveform_sig_loopback =1672;
31533: waveform_sig_loopback =-340;
31534: waveform_sig_loopback =1241;
31535: waveform_sig_loopback =-243;
31536: waveform_sig_loopback =449;
31537: waveform_sig_loopback =1787;
31538: waveform_sig_loopback =-532;
31539: waveform_sig_loopback =1049;
31540: waveform_sig_loopback =918;
31541: waveform_sig_loopback =772;
31542: waveform_sig_loopback =99;
31543: waveform_sig_loopback =2059;
31544: waveform_sig_loopback =472;
31545: waveform_sig_loopback =209;
31546: waveform_sig_loopback =2136;
31547: waveform_sig_loopback =658;
31548: waveform_sig_loopback =737;
31549: waveform_sig_loopback =1321;
31550: waveform_sig_loopback =1951;
31551: waveform_sig_loopback =365;
31552: waveform_sig_loopback =906;
31553: waveform_sig_loopback =2812;
31554: waveform_sig_loopback =686;
31555: waveform_sig_loopback =196;
31556: waveform_sig_loopback =3005;
31557: waveform_sig_loopback =1892;
31558: waveform_sig_loopback =-78;
31559: waveform_sig_loopback =2124;
31560: waveform_sig_loopback =2945;
31561: waveform_sig_loopback =235;
31562: waveform_sig_loopback =3712;
31563: waveform_sig_loopback =127;
31564: waveform_sig_loopback =-53;
31565: waveform_sig_loopback =4900;
31566: waveform_sig_loopback =1603;
31567: waveform_sig_loopback =1455;
31568: waveform_sig_loopback =753;
31569: waveform_sig_loopback =2533;
31570: waveform_sig_loopback =4031;
31571: waveform_sig_loopback =929;
31572: waveform_sig_loopback =1461;
31573: waveform_sig_loopback =3161;
31574: waveform_sig_loopback =1642;
31575: waveform_sig_loopback =3295;
31576: waveform_sig_loopback =1182;
31577: waveform_sig_loopback =2627;
31578: waveform_sig_loopback =3521;
31579: waveform_sig_loopback =1188;
31580: waveform_sig_loopback =3141;
31581: waveform_sig_loopback =2558;
31582: waveform_sig_loopback =2553;
31583: waveform_sig_loopback =2163;
31584: waveform_sig_loopback =3728;
31585: waveform_sig_loopback =2200;
31586: waveform_sig_loopback =2289;
31587: waveform_sig_loopback =3699;
31588: waveform_sig_loopback =2654;
31589: waveform_sig_loopback =2524;
31590: waveform_sig_loopback =2934;
31591: waveform_sig_loopback =4109;
31592: waveform_sig_loopback =1804;
31593: waveform_sig_loopback =2851;
31594: waveform_sig_loopback =4801;
31595: waveform_sig_loopback =2017;
31596: waveform_sig_loopback =2373;
31597: waveform_sig_loopback =4689;
31598: waveform_sig_loopback =3413;
31599: waveform_sig_loopback =1987;
31600: waveform_sig_loopback =3751;
31601: waveform_sig_loopback =4668;
31602: waveform_sig_loopback =2163;
31603: waveform_sig_loopback =5304;
31604: waveform_sig_loopback =1787;
31605: waveform_sig_loopback =1969;
31606: waveform_sig_loopback =6424;
31607: waveform_sig_loopback =3533;
31608: waveform_sig_loopback =2956;
31609: waveform_sig_loopback =2504;
31610: waveform_sig_loopback =4592;
31611: waveform_sig_loopback =5330;
31612: waveform_sig_loopback =2761;
31613: waveform_sig_loopback =3311;
31614: waveform_sig_loopback =4609;
31615: waveform_sig_loopback =3569;
31616: waveform_sig_loopback =4801;
31617: waveform_sig_loopback =2866;
31618: waveform_sig_loopback =4570;
31619: waveform_sig_loopback =4883;
31620: waveform_sig_loopback =2986;
31621: waveform_sig_loopback =4828;
31622: waveform_sig_loopback =4068;
31623: waveform_sig_loopback =4269;
31624: waveform_sig_loopback =3853;
31625: waveform_sig_loopback =5224;
31626: waveform_sig_loopback =3936;
31627: waveform_sig_loopback =3877;
31628: waveform_sig_loopback =5167;
31629: waveform_sig_loopback =4563;
31630: waveform_sig_loopback =3696;
31631: waveform_sig_loopback =4819;
31632: waveform_sig_loopback =5715;
31633: waveform_sig_loopback =2968;
31634: waveform_sig_loopback =4993;
31635: waveform_sig_loopback =6035;
31636: waveform_sig_loopback =3518;
31637: waveform_sig_loopback =4313;
31638: waveform_sig_loopback =5891;
31639: waveform_sig_loopback =5196;
31640: waveform_sig_loopback =3475;
31641: waveform_sig_loopback =5184;
31642: waveform_sig_loopback =6438;
31643: waveform_sig_loopback =3408;
31644: waveform_sig_loopback =6982;
31645: waveform_sig_loopback =3147;
31646: waveform_sig_loopback =3470;
31647: waveform_sig_loopback =8127;
31648: waveform_sig_loopback =4781;
31649: waveform_sig_loopback =4342;
31650: waveform_sig_loopback =4185;
31651: waveform_sig_loopback =6029;
31652: waveform_sig_loopback =6638;
31653: waveform_sig_loopback =4249;
31654: waveform_sig_loopback =4846;
31655: waveform_sig_loopback =5969;
31656: waveform_sig_loopback =5155;
31657: waveform_sig_loopback =5997;
31658: waveform_sig_loopback =4363;
31659: waveform_sig_loopback =6197;
31660: waveform_sig_loopback =5892;
31661: waveform_sig_loopback =4685;
31662: waveform_sig_loopback =6142;
31663: waveform_sig_loopback =5300;
31664: waveform_sig_loopback =5947;
31665: waveform_sig_loopback =4819;
31666: waveform_sig_loopback =6768;
31667: waveform_sig_loopback =5340;
31668: waveform_sig_loopback =4878;
31669: waveform_sig_loopback =6947;
31670: waveform_sig_loopback =5506;
31671: waveform_sig_loopback =5002;
31672: waveform_sig_loopback =6538;
31673: waveform_sig_loopback =6395;
31674: waveform_sig_loopback =4636;
31675: waveform_sig_loopback =6256;
31676: waveform_sig_loopback =7058;
31677: waveform_sig_loopback =4963;
31678: waveform_sig_loopback =5361;
31679: waveform_sig_loopback =7245;
31680: waveform_sig_loopback =6308;
31681: waveform_sig_loopback =4594;
31682: waveform_sig_loopback =6572;
31683: waveform_sig_loopback =7500;
31684: waveform_sig_loopback =4535;
31685: waveform_sig_loopback =8218;
31686: waveform_sig_loopback =4206;
31687: waveform_sig_loopback =4709;
31688: waveform_sig_loopback =9355;
31689: waveform_sig_loopback =5822;
31690: waveform_sig_loopback =5338;
31691: waveform_sig_loopback =5542;
31692: waveform_sig_loopback =7014;
31693: waveform_sig_loopback =7788;
31694: waveform_sig_loopback =5413;
31695: waveform_sig_loopback =5646;
31696: waveform_sig_loopback =7270;
31697: waveform_sig_loopback =6172;
31698: waveform_sig_loopback =6805;
31699: waveform_sig_loopback =5690;
31700: waveform_sig_loopback =6982;
31701: waveform_sig_loopback =6957;
31702: waveform_sig_loopback =5900;
31703: waveform_sig_loopback =6704;
31704: waveform_sig_loopback =6687;
31705: waveform_sig_loopback =6720;
31706: waveform_sig_loopback =5704;
31707: waveform_sig_loopback =8141;
31708: waveform_sig_loopback =5704;
31709: waveform_sig_loopback =6191;
31710: waveform_sig_loopback =7872;
31711: waveform_sig_loopback =6176;
31712: waveform_sig_loopback =6247;
31713: waveform_sig_loopback =7246;
31714: waveform_sig_loopback =7306;
31715: waveform_sig_loopback =5558;
31716: waveform_sig_loopback =7084;
31717: waveform_sig_loopback =7899;
31718: waveform_sig_loopback =5773;
31719: waveform_sig_loopback =6238;
31720: waveform_sig_loopback =8073;
31721: waveform_sig_loopback =7113;
31722: waveform_sig_loopback =5228;
31723: waveform_sig_loopback =7593;
31724: waveform_sig_loopback =8209;
31725: waveform_sig_loopback =5162;
31726: waveform_sig_loopback =9308;
31727: waveform_sig_loopback =4507;
31728: waveform_sig_loopback =5650;
31729: waveform_sig_loopback =10317;
31730: waveform_sig_loopback =6026;
31731: waveform_sig_loopback =6298;
31732: waveform_sig_loopback =6219;
31733: waveform_sig_loopback =7449;
31734: waveform_sig_loopback =8862;
31735: waveform_sig_loopback =5608;
31736: waveform_sig_loopback =6483;
31737: waveform_sig_loopback =8083;
31738: waveform_sig_loopback =6339;
31739: waveform_sig_loopback =7850;
31740: waveform_sig_loopback =6040;
31741: waveform_sig_loopback =7480;
31742: waveform_sig_loopback =7829;
31743: waveform_sig_loopback =6053;
31744: waveform_sig_loopback =7517;
31745: waveform_sig_loopback =7319;
31746: waveform_sig_loopback =6917;
31747: waveform_sig_loopback =6637;
31748: waveform_sig_loopback =8367;
31749: waveform_sig_loopback =6253;
31750: waveform_sig_loopback =6911;
31751: waveform_sig_loopback =8097;
31752: waveform_sig_loopback =6747;
31753: waveform_sig_loopback =6636;
31754: waveform_sig_loopback =7816;
31755: waveform_sig_loopback =7566;
31756: waveform_sig_loopback =6065;
31757: waveform_sig_loopback =7537;
31758: waveform_sig_loopback =8224;
31759: waveform_sig_loopback =6296;
31760: waveform_sig_loopback =6333;
31761: waveform_sig_loopback =8824;
31762: waveform_sig_loopback =7238;
31763: waveform_sig_loopback =5376;
31764: waveform_sig_loopback =8504;
31765: waveform_sig_loopback =7828;
31766: waveform_sig_loopback =5924;
31767: waveform_sig_loopback =9601;
31768: waveform_sig_loopback =4197;
31769: waveform_sig_loopback =6850;
31770: waveform_sig_loopback =9944;
31771: waveform_sig_loopback =6443;
31772: waveform_sig_loopback =6794;
31773: waveform_sig_loopback =5963;
31774: waveform_sig_loopback =8237;
31775: waveform_sig_loopback =8790;
31776: waveform_sig_loopback =5632;
31777: waveform_sig_loopback =7165;
31778: waveform_sig_loopback =7813;
31779: waveform_sig_loopback =6777;
31780: waveform_sig_loopback =8056;
31781: waveform_sig_loopback =5944;
31782: waveform_sig_loopback =8010;
31783: waveform_sig_loopback =7688;
31784: waveform_sig_loopback =6163;
31785: waveform_sig_loopback =7780;
31786: waveform_sig_loopback =7232;
31787: waveform_sig_loopback =7000;
31788: waveform_sig_loopback =6780;
31789: waveform_sig_loopback =8375;
31790: waveform_sig_loopback =6137;
31791: waveform_sig_loopback =7189;
31792: waveform_sig_loopback =7904;
31793: waveform_sig_loopback =6740;
31794: waveform_sig_loopback =6773;
31795: waveform_sig_loopback =7538;
31796: waveform_sig_loopback =7789;
31797: waveform_sig_loopback =5804;
31798: waveform_sig_loopback =7467;
31799: waveform_sig_loopback =8453;
31800: waveform_sig_loopback =5719;
31801: waveform_sig_loopback =6623;
31802: waveform_sig_loopback =8752;
31803: waveform_sig_loopback =6705;
31804: waveform_sig_loopback =5707;
31805: waveform_sig_loopback =8157;
31806: waveform_sig_loopback =7544;
31807: waveform_sig_loopback =6102;
31808: waveform_sig_loopback =8977;
31809: waveform_sig_loopback =4132;
31810: waveform_sig_loopback =6871;
31811: waveform_sig_loopback =9410;
31812: waveform_sig_loopback =6518;
31813: waveform_sig_loopback =6212;
31814: waveform_sig_loopback =5815;
31815: waveform_sig_loopback =8229;
31816: waveform_sig_loopback =8099;
31817: waveform_sig_loopback =5469;
31818: waveform_sig_loopback =6844;
31819: waveform_sig_loopback =7324;
31820: waveform_sig_loopback =6644;
31821: waveform_sig_loopback =7578;
31822: waveform_sig_loopback =5448;
31823: waveform_sig_loopback =7869;
31824: waveform_sig_loopback =7082;
31825: waveform_sig_loopback =5844;
31826: waveform_sig_loopback =7474;
31827: waveform_sig_loopback =6598;
31828: waveform_sig_loopback =6623;
31829: waveform_sig_loopback =6484;
31830: waveform_sig_loopback =7624;
31831: waveform_sig_loopback =5860;
31832: waveform_sig_loopback =6475;
31833: waveform_sig_loopback =7290;
31834: waveform_sig_loopback =6657;
31835: waveform_sig_loopback =5825;
31836: waveform_sig_loopback =7141;
31837: waveform_sig_loopback =7166;
31838: waveform_sig_loopback =5107;
31839: waveform_sig_loopback =7335;
31840: waveform_sig_loopback =7413;
31841: waveform_sig_loopback =5007;
31842: waveform_sig_loopback =6533;
31843: waveform_sig_loopback =7792;
31844: waveform_sig_loopback =6064;
31845: waveform_sig_loopback =5135;
31846: waveform_sig_loopback =7404;
31847: waveform_sig_loopback =7072;
31848: waveform_sig_loopback =5222;
31849: waveform_sig_loopback =8257;
31850: waveform_sig_loopback =3568;
31851: waveform_sig_loopback =6063;
31852: waveform_sig_loopback =8738;
31853: waveform_sig_loopback =5718;
31854: waveform_sig_loopback =5261;
31855: waveform_sig_loopback =5348;
31856: waveform_sig_loopback =7303;
31857: waveform_sig_loopback =7183;
31858: waveform_sig_loopback =4812;
31859: waveform_sig_loopback =5984;
31860: waveform_sig_loopback =6451;
31861: waveform_sig_loopback =5931;
31862: waveform_sig_loopback =6504;
31863: waveform_sig_loopback =4740;
31864: waveform_sig_loopback =7110;
31865: waveform_sig_loopback =5873;
31866: waveform_sig_loopback =5265;
31867: waveform_sig_loopback =6475;
31868: waveform_sig_loopback =5571;
31869: waveform_sig_loopback =5988;
31870: waveform_sig_loopback =5306;
31871: waveform_sig_loopback =6847;
31872: waveform_sig_loopback =4911;
31873: waveform_sig_loopback =5448;
31874: waveform_sig_loopback =6641;
31875: waveform_sig_loopback =5309;
31876: waveform_sig_loopback =4854;
31877: waveform_sig_loopback =6626;
31878: waveform_sig_loopback =5787;
31879: waveform_sig_loopback =4150;
31880: waveform_sig_loopback =6436;
31881: waveform_sig_loopback =6218;
31882: waveform_sig_loopback =4176;
31883: waveform_sig_loopback =5296;
31884: waveform_sig_loopback =6653;
31885: waveform_sig_loopback =5162;
31886: waveform_sig_loopback =3981;
31887: waveform_sig_loopback =6317;
31888: waveform_sig_loopback =5974;
31889: waveform_sig_loopback =4070;
31890: waveform_sig_loopback =7219;
31891: waveform_sig_loopback =2262;
31892: waveform_sig_loopback =4959;
31893: waveform_sig_loopback =7874;
31894: waveform_sig_loopback =4274;
31895: waveform_sig_loopback =3980;
31896: waveform_sig_loopback =4527;
31897: waveform_sig_loopback =5926;
31898: waveform_sig_loopback =6104;
31899: waveform_sig_loopback =3546;
31900: waveform_sig_loopback =4704;
31901: waveform_sig_loopback =5499;
31902: waveform_sig_loopback =4528;
31903: waveform_sig_loopback =5177;
31904: waveform_sig_loopback =3725;
31905: waveform_sig_loopback =5708;
31906: waveform_sig_loopback =4593;
31907: waveform_sig_loopback =4091;
31908: waveform_sig_loopback =5024;
31909: waveform_sig_loopback =4457;
31910: waveform_sig_loopback =4555;
31911: waveform_sig_loopback =3897;
31912: waveform_sig_loopback =5763;
31913: waveform_sig_loopback =3360;
31914: waveform_sig_loopback =4116;
31915: waveform_sig_loopback =5475;
31916: waveform_sig_loopback =3633;
31917: waveform_sig_loopback =3712;
31918: waveform_sig_loopback =5308;
31919: waveform_sig_loopback =4054;
31920: waveform_sig_loopback =3149;
31921: waveform_sig_loopback =4903;
31922: waveform_sig_loopback =4668;
31923: waveform_sig_loopback =3019;
31924: waveform_sig_loopback =3632;
31925: waveform_sig_loopback =5469;
31926: waveform_sig_loopback =3580;
31927: waveform_sig_loopback =2317;
31928: waveform_sig_loopback =5400;
31929: waveform_sig_loopback =4060;
31930: waveform_sig_loopback =2758;
31931: waveform_sig_loopback =5857;
31932: waveform_sig_loopback =396;
31933: waveform_sig_loopback =3968;
31934: waveform_sig_loopback =6157;
31935: waveform_sig_loopback =2569;
31936: waveform_sig_loopback =2693;
31937: waveform_sig_loopback =2955;
31938: waveform_sig_loopback =4388;
31939: waveform_sig_loopback =4729;
31940: waveform_sig_loopback =1746;
31941: waveform_sig_loopback =3308;
31942: waveform_sig_loopback =4004;
31943: waveform_sig_loopback =2772;
31944: waveform_sig_loopback =3816;
31945: waveform_sig_loopback =2087;
31946: waveform_sig_loopback =4053;
31947: waveform_sig_loopback =3143;
31948: waveform_sig_loopback =2406;
31949: waveform_sig_loopback =3343;
31950: waveform_sig_loopback =3087;
31951: waveform_sig_loopback =2647;
31952: waveform_sig_loopback =2505;
31953: waveform_sig_loopback =4181;
31954: waveform_sig_loopback =1366;
31955: waveform_sig_loopback =2972;
31956: waveform_sig_loopback =3567;
31957: waveform_sig_loopback =1824;
31958: waveform_sig_loopback =2383;
31959: waveform_sig_loopback =3295;
31960: waveform_sig_loopback =2469;
31961: waveform_sig_loopback =1543;
31962: waveform_sig_loopback =3002;
31963: waveform_sig_loopback =3253;
31964: waveform_sig_loopback =1063;
31965: waveform_sig_loopback =1990;
31966: waveform_sig_loopback =4002;
31967: waveform_sig_loopback =1543;
31968: waveform_sig_loopback =789;
31969: waveform_sig_loopback =3784;
31970: waveform_sig_loopback =1971;
31971: waveform_sig_loopback =1433;
31972: waveform_sig_loopback =3949;
31973: waveform_sig_loopback =-1605;
31974: waveform_sig_loopback =2708;
31975: waveform_sig_loopback =4075;
31976: waveform_sig_loopback =836;
31977: waveform_sig_loopback =1087;
31978: waveform_sig_loopback =948;
31979: waveform_sig_loopback =2869;
31980: waveform_sig_loopback =2839;
31981: waveform_sig_loopback =-326;
31982: waveform_sig_loopback =1849;
31983: waveform_sig_loopback =1977;
31984: waveform_sig_loopback =933;
31985: waveform_sig_loopback =2195;
31986: waveform_sig_loopback =-9;
31987: waveform_sig_loopback =2486;
31988: waveform_sig_loopback =1288;
31989: waveform_sig_loopback =369;
31990: waveform_sig_loopback =1749;
31991: waveform_sig_loopback =1108;
31992: waveform_sig_loopback =648;
31993: waveform_sig_loopback =1090;
31994: waveform_sig_loopback =1935;
31995: waveform_sig_loopback =-389;
31996: waveform_sig_loopback =1362;
31997: waveform_sig_loopback =1349;
31998: waveform_sig_loopback =334;
31999: waveform_sig_loopback =360;
32000: waveform_sig_loopback =1499;
32001: waveform_sig_loopback =848;
32002: waveform_sig_loopback =-621;
32003: waveform_sig_loopback =1408;
32004: waveform_sig_loopback =1337;
32005: waveform_sig_loopback =-961;
32006: waveform_sig_loopback =417;
32007: waveform_sig_loopback =1965;
32008: waveform_sig_loopback =-404;
32009: waveform_sig_loopback =-880;
32010: waveform_sig_loopback =1919;
32011: waveform_sig_loopback =-127;
32012: waveform_sig_loopback =-165;
32013: waveform_sig_loopback =1854;
32014: waveform_sig_loopback =-3561;
32015: waveform_sig_loopback =1288;
32016: waveform_sig_loopback =1827;
32017: waveform_sig_loopback =-892;
32018: waveform_sig_loopback =-825;
32019: waveform_sig_loopback =-1143;
32020: waveform_sig_loopback =1464;
32021: waveform_sig_loopback =556;
32022: waveform_sig_loopback =-2139;
32023: waveform_sig_loopback =336;
32024: waveform_sig_loopback =-407;
32025: waveform_sig_loopback =-392;
32026: waveform_sig_loopback =-32;
32027: waveform_sig_loopback =-1934;
32028: waveform_sig_loopback =1008;
32029: waveform_sig_loopback =-1075;
32030: waveform_sig_loopback =-1212;
32031: waveform_sig_loopback =-128;
32032: waveform_sig_loopback =-942;
32033: waveform_sig_loopback =-1016;
32034: waveform_sig_loopback =-918;
32035: waveform_sig_loopback =-2;
32036: waveform_sig_loopback =-2154;
32037: waveform_sig_loopback =-563;
32038: waveform_sig_loopback =-563;
32039: waveform_sig_loopback =-1500;
32040: waveform_sig_loopback =-1568;
32041: waveform_sig_loopback =-390;
32042: waveform_sig_loopback =-1075;
32043: waveform_sig_loopback =-2670;
32044: waveform_sig_loopback =-243;
32045: waveform_sig_loopback =-625;
32046: waveform_sig_loopback =-3128;
32047: waveform_sig_loopback =-1022;
32048: waveform_sig_loopback =-200;
32049: waveform_sig_loopback =-2413;
32050: waveform_sig_loopback =-2487;
32051: waveform_sig_loopback =-285;
32052: waveform_sig_loopback =-1787;
32053: waveform_sig_loopback =-2012;
32054: waveform_sig_loopback =-346;
32055: waveform_sig_loopback =-5185;
32056: waveform_sig_loopback =-669;
32057: waveform_sig_loopback =-54;
32058: waveform_sig_loopback =-2665;
32059: waveform_sig_loopback =-2966;
32060: waveform_sig_loopback =-2662;
32061: waveform_sig_loopback =-445;
32062: waveform_sig_loopback =-1586;
32063: waveform_sig_loopback =-3721;
32064: waveform_sig_loopback =-1681;
32065: waveform_sig_loopback =-2313;
32066: waveform_sig_loopback =-2037;
32067: waveform_sig_loopback =-2241;
32068: waveform_sig_loopback =-3500;
32069: waveform_sig_loopback =-923;
32070: waveform_sig_loopback =-3164;
32071: waveform_sig_loopback =-2731;
32072: waveform_sig_loopback =-2208;
32073: waveform_sig_loopback =-2748;
32074: waveform_sig_loopback =-2837;
32075: waveform_sig_loopback =-2802;
32076: waveform_sig_loopback =-1847;
32077: waveform_sig_loopback =-3950;
32078: waveform_sig_loopback =-2448;
32079: waveform_sig_loopback =-2320;
32080: waveform_sig_loopback =-3305;
32081: waveform_sig_loopback =-3552;
32082: waveform_sig_loopback =-1873;
32083: waveform_sig_loopback =-3162;
32084: waveform_sig_loopback =-4466;
32085: waveform_sig_loopback =-1722;
32086: waveform_sig_loopback =-2931;
32087: waveform_sig_loopback =-4644;
32088: waveform_sig_loopback =-2719;
32089: waveform_sig_loopback =-2314;
32090: waveform_sig_loopback =-3857;
32091: waveform_sig_loopback =-4531;
32092: waveform_sig_loopback =-1918;
32093: waveform_sig_loopback =-3521;
32094: waveform_sig_loopback =-3985;
32095: waveform_sig_loopback =-1889;
32096: waveform_sig_loopback =-7110;
32097: waveform_sig_loopback =-2287;
32098: waveform_sig_loopback =-1677;
32099: waveform_sig_loopback =-4749;
32100: waveform_sig_loopback =-4603;
32101: waveform_sig_loopback =-4215;
32102: waveform_sig_loopback =-2406;
32103: waveform_sig_loopback =-3194;
32104: waveform_sig_loopback =-5463;
32105: waveform_sig_loopback =-3403;
32106: waveform_sig_loopback =-3897;
32107: waveform_sig_loopback =-3820;
32108: waveform_sig_loopback =-4027;
32109: waveform_sig_loopback =-4954;
32110: waveform_sig_loopback =-2726;
32111: waveform_sig_loopback =-4873;
32112: waveform_sig_loopback =-4242;
32113: waveform_sig_loopback =-4058;
32114: waveform_sig_loopback =-4214;
32115: waveform_sig_loopback =-4484;
32116: waveform_sig_loopback =-4582;
32117: waveform_sig_loopback =-3245;
32118: waveform_sig_loopback =-5755;
32119: waveform_sig_loopback =-4121;
32120: waveform_sig_loopback =-3655;
32121: waveform_sig_loopback =-5341;
32122: waveform_sig_loopback =-4796;
32123: waveform_sig_loopback =-3443;
32124: waveform_sig_loopback =-5167;
32125: waveform_sig_loopback =-5471;
32126: waveform_sig_loopback =-3562;
32127: waveform_sig_loopback =-4481;
32128: waveform_sig_loopback =-6060;
32129: waveform_sig_loopback =-4545;
32130: waveform_sig_loopback =-3492;
32131: waveform_sig_loopback =-5587;
32132: waveform_sig_loopback =-6085;
32133: waveform_sig_loopback =-3104;
32134: waveform_sig_loopback =-5405;
32135: waveform_sig_loopback =-5171;
32136: waveform_sig_loopback =-3562;
32137: waveform_sig_loopback =-8688;
32138: waveform_sig_loopback =-3467;
32139: waveform_sig_loopback =-3312;
32140: waveform_sig_loopback =-6223;
32141: waveform_sig_loopback =-6062;
32142: waveform_sig_loopback =-5522;
32143: waveform_sig_loopback =-3927;
32144: waveform_sig_loopback =-4635;
32145: waveform_sig_loopback =-6921;
32146: waveform_sig_loopback =-4866;
32147: waveform_sig_loopback =-5109;
32148: waveform_sig_loopback =-5445;
32149: waveform_sig_loopback =-5385;
32150: waveform_sig_loopback =-6168;
32151: waveform_sig_loopback =-4429;
32152: waveform_sig_loopback =-5934;
32153: waveform_sig_loopback =-5736;
32154: waveform_sig_loopback =-5511;
32155: waveform_sig_loopback =-5196;
32156: waveform_sig_loopback =-6335;
32157: waveform_sig_loopback =-5509;
32158: waveform_sig_loopback =-4653;
32159: waveform_sig_loopback =-7419;
32160: waveform_sig_loopback =-4900;
32161: waveform_sig_loopback =-5400;
32162: waveform_sig_loopback =-6493;
32163: waveform_sig_loopback =-6002;
32164: waveform_sig_loopback =-5004;
32165: waveform_sig_loopback =-6201;
32166: waveform_sig_loopback =-6881;
32167: waveform_sig_loopback =-4805;
32168: waveform_sig_loopback =-5758;
32169: waveform_sig_loopback =-7337;
32170: waveform_sig_loopback =-5689;
32171: waveform_sig_loopback =-4718;
32172: waveform_sig_loopback =-6989;
32173: waveform_sig_loopback =-7286;
32174: waveform_sig_loopback =-4065;
32175: waveform_sig_loopback =-6917;
32176: waveform_sig_loopback =-6124;
32177: waveform_sig_loopback =-4774;
32178: waveform_sig_loopback =-10152;
32179: waveform_sig_loopback =-4054;
32180: waveform_sig_loopback =-4846;
32181: waveform_sig_loopback =-7488;
32182: waveform_sig_loopback =-7008;
32183: waveform_sig_loopback =-6972;
32184: waveform_sig_loopback =-4641;
32185: waveform_sig_loopback =-5798;
32186: waveform_sig_loopback =-8509;
32187: waveform_sig_loopback =-5582;
32188: waveform_sig_loopback =-6262;
32189: waveform_sig_loopback =-6533;
32190: waveform_sig_loopback =-6278;
32191: waveform_sig_loopback =-7620;
32192: waveform_sig_loopback =-5078;
32193: waveform_sig_loopback =-6975;
32194: waveform_sig_loopback =-7136;
32195: waveform_sig_loopback =-6136;
32196: waveform_sig_loopback =-6435;
32197: waveform_sig_loopback =-7334;
32198: waveform_sig_loopback =-6200;
32199: waveform_sig_loopback =-6072;
32200: waveform_sig_loopback =-7942;
32201: waveform_sig_loopback =-5855;
32202: waveform_sig_loopback =-6578;
32203: waveform_sig_loopback =-7247;
32204: waveform_sig_loopback =-6885;
32205: waveform_sig_loopback =-5861;
32206: waveform_sig_loopback =-7221;
32207: waveform_sig_loopback =-7700;
32208: waveform_sig_loopback =-5611;
32209: waveform_sig_loopback =-6579;
32210: waveform_sig_loopback =-8284;
32211: waveform_sig_loopback =-6455;
32212: waveform_sig_loopback =-5345;
32213: waveform_sig_loopback =-8155;
32214: waveform_sig_loopback =-7816;
32215: waveform_sig_loopback =-4837;
32216: waveform_sig_loopback =-8097;
32217: waveform_sig_loopback =-6301;
32218: waveform_sig_loopback =-6129;
32219: waveform_sig_loopback =-10746;
32220: waveform_sig_loopback =-4315;
32221: waveform_sig_loopback =-6202;
32222: waveform_sig_loopback =-7772;
32223: waveform_sig_loopback =-7692;
32224: waveform_sig_loopback =-7753;
32225: waveform_sig_loopback =-4911;
32226: waveform_sig_loopback =-7035;
32227: waveform_sig_loopback =-8739;
32228: waveform_sig_loopback =-5931;
32229: waveform_sig_loopback =-7592;
32230: waveform_sig_loopback =-6549;
32231: waveform_sig_loopback =-7293;
32232: waveform_sig_loopback =-8047;
32233: waveform_sig_loopback =-5493;
32234: waveform_sig_loopback =-8137;
32235: waveform_sig_loopback =-7137;
32236: waveform_sig_loopback =-6926;
32237: waveform_sig_loopback =-6996;
32238: waveform_sig_loopback =-7806;
32239: waveform_sig_loopback =-6709;
32240: waveform_sig_loopback =-6581;
32241: waveform_sig_loopback =-8595;
32242: waveform_sig_loopback =-6111;
32243: waveform_sig_loopback =-7299;
32244: waveform_sig_loopback =-7466;
32245: waveform_sig_loopback =-7473;
32246: waveform_sig_loopback =-6409;
32247: waveform_sig_loopback =-7320;
32248: waveform_sig_loopback =-8500;
32249: waveform_sig_loopback =-5657;
32250: waveform_sig_loopback =-7144;
32251: waveform_sig_loopback =-8908;
32252: waveform_sig_loopback =-6215;
32253: waveform_sig_loopback =-6270;
32254: waveform_sig_loopback =-8356;
32255: waveform_sig_loopback =-7801;
32256: waveform_sig_loopback =-5557;
32257: waveform_sig_loopback =-8107;
32258: waveform_sig_loopback =-6594;
32259: waveform_sig_loopback =-6784;
32260: waveform_sig_loopback =-10539;
32261: waveform_sig_loopback =-4872;
32262: waveform_sig_loopback =-6372;
32263: waveform_sig_loopback =-7885;
32264: waveform_sig_loopback =-8353;
32265: waveform_sig_loopback =-7506;
32266: waveform_sig_loopback =-5307;
32267: waveform_sig_loopback =-7371;
32268: waveform_sig_loopback =-8614;
32269: waveform_sig_loopback =-6341;
32270: waveform_sig_loopback =-7613;
32271: waveform_sig_loopback =-6580;
32272: waveform_sig_loopback =-7575;
32273: waveform_sig_loopback =-7947;
32274: waveform_sig_loopback =-5637;
32275: waveform_sig_loopback =-8268;
32276: waveform_sig_loopback =-7073;
32277: waveform_sig_loopback =-6971;
32278: waveform_sig_loopback =-7251;
32279: waveform_sig_loopback =-7624;
32280: waveform_sig_loopback =-6767;
32281: waveform_sig_loopback =-6803;
32282: waveform_sig_loopback =-8258;
32283: waveform_sig_loopback =-6463;
32284: waveform_sig_loopback =-7001;
32285: waveform_sig_loopback =-7491;
32286: waveform_sig_loopback =-7667;
32287: waveform_sig_loopback =-5894;
32288: waveform_sig_loopback =-7721;
32289: waveform_sig_loopback =-8227;
32290: waveform_sig_loopback =-5399;
32291: waveform_sig_loopback =-7482;
32292: waveform_sig_loopback =-8414;
32293: waveform_sig_loopback =-6158;
32294: waveform_sig_loopback =-6323;
32295: waveform_sig_loopback =-8006;
32296: waveform_sig_loopback =-7773;
32297: waveform_sig_loopback =-5339;
32298: waveform_sig_loopback =-7864;
32299: waveform_sig_loopback =-6490;
32300: waveform_sig_loopback =-6573;
32301: waveform_sig_loopback =-10243;
32302: waveform_sig_loopback =-4658;
32303: waveform_sig_loopback =-5974;
32304: waveform_sig_loopback =-7873;
32305: waveform_sig_loopback =-8030;
32306: waveform_sig_loopback =-6909;
32307: waveform_sig_loopback =-5337;
32308: waveform_sig_loopback =-6964;
32309: waveform_sig_loopback =-8248;
32310: waveform_sig_loopback =-6149;
32311: waveform_sig_loopback =-7100;
32312: waveform_sig_loopback =-6424;
32313: waveform_sig_loopback =-7221;
32314: waveform_sig_loopback =-7351;
32315: waveform_sig_loopback =-5468;
32316: waveform_sig_loopback =-7852;
32317: waveform_sig_loopback =-6527;
32318: waveform_sig_loopback =-6631;
32319: waveform_sig_loopback =-6817;
32320: waveform_sig_loopback =-7046;
32321: waveform_sig_loopback =-6465;
32322: waveform_sig_loopback =-6141;
32323: waveform_sig_loopback =-7850;
32324: waveform_sig_loopback =-6136;
32325: waveform_sig_loopback =-6062;
32326: waveform_sig_loopback =-7480;
32327: waveform_sig_loopback =-6725;
32328: waveform_sig_loopback =-5326;
32329: waveform_sig_loopback =-7589;
32330: waveform_sig_loopback =-7020;
32331: waveform_sig_loopback =-5235;
32332: waveform_sig_loopback =-6827;
32333: waveform_sig_loopback =-7598;
32334: waveform_sig_loopback =-5807;
32335: waveform_sig_loopback =-5469;
32336: waveform_sig_loopback =-7569;
32337: waveform_sig_loopback =-7069;
32338: waveform_sig_loopback =-4478;
32339: waveform_sig_loopback =-7460;
32340: waveform_sig_loopback =-5605;
32341: waveform_sig_loopback =-5976;
32342: waveform_sig_loopback =-9552;
32343: waveform_sig_loopback =-3750;
32344: waveform_sig_loopback =-5333;
32345: waveform_sig_loopback =-7283;
32346: waveform_sig_loopback =-7150;
32347: waveform_sig_loopback =-6104;
32348: waveform_sig_loopback =-4728;
32349: waveform_sig_loopback =-6066;
32350: waveform_sig_loopback =-7586;
32351: waveform_sig_loopback =-5303;
32352: waveform_sig_loopback =-6117;
32353: waveform_sig_loopback =-5803;
32354: waveform_sig_loopback =-6314;
32355: waveform_sig_loopback =-6414;
32356: waveform_sig_loopback =-4800;
32357: waveform_sig_loopback =-6785;
32358: waveform_sig_loopback =-5771;
32359: waveform_sig_loopback =-5833;
32360: waveform_sig_loopback =-5675;
32361: waveform_sig_loopback =-6438;
32362: waveform_sig_loopback =-5337;
32363: waveform_sig_loopback =-5228;
32364: waveform_sig_loopback =-7110;
32365: waveform_sig_loopback =-4827;
32366: waveform_sig_loopback =-5278;
32367: waveform_sig_loopback =-6679;
32368: waveform_sig_loopback =-5362;
32369: waveform_sig_loopback =-4655;
32370: waveform_sig_loopback =-6562;
32371: waveform_sig_loopback =-5762;
32372: waveform_sig_loopback =-4477;
32373: waveform_sig_loopback =-5592;
32374: waveform_sig_loopback =-6664;
32375: waveform_sig_loopback =-4775;
32376: waveform_sig_loopback =-4198;
32377: waveform_sig_loopback =-6826;
32378: waveform_sig_loopback =-5725;
32379: waveform_sig_loopback =-3328;
32380: waveform_sig_loopback =-6700;
32381: waveform_sig_loopback =-4079;
32382: waveform_sig_loopback =-5270;
32383: waveform_sig_loopback =-8372;
32384: waveform_sig_loopback =-2306;
32385: waveform_sig_loopback =-4522;
32386: waveform_sig_loopback =-6078;
32387: waveform_sig_loopback =-5884;
32388: waveform_sig_loopback =-5008;
32389: waveform_sig_loopback =-3341;
32390: waveform_sig_loopback =-4981;
32391: waveform_sig_loopback =-6458;
32392: waveform_sig_loopback =-3850;
32393: waveform_sig_loopback =-5035;
32394: waveform_sig_loopback =-4566;
32395: waveform_sig_loopback =-5011;
32396: waveform_sig_loopback =-5217;
32397: waveform_sig_loopback =-3516;
32398: waveform_sig_loopback =-5401;
32399: waveform_sig_loopback =-4641;
32400: waveform_sig_loopback =-4417;
32401: waveform_sig_loopback =-4296;
32402: waveform_sig_loopback =-5404;
32403: waveform_sig_loopback =-3570;
32404: waveform_sig_loopback =-4252;
32405: waveform_sig_loopback =-5691;
32406: waveform_sig_loopback =-3145;
32407: waveform_sig_loopback =-4468;
32408: waveform_sig_loopback =-4897;
32409: waveform_sig_loopback =-4093;
32410: waveform_sig_loopback =-3464;
32411: waveform_sig_loopback =-4817;
32412: waveform_sig_loopback =-4707;
32413: waveform_sig_loopback =-2868;
32414: waveform_sig_loopback =-4203;
32415: waveform_sig_loopback =-5447;
32416: waveform_sig_loopback =-2974;
32417: waveform_sig_loopback =-2986;
32418: waveform_sig_loopback =-5453;
32419: waveform_sig_loopback =-4001;
32420: waveform_sig_loopback =-2068;
32421: waveform_sig_loopback =-5225;
32422: waveform_sig_loopback =-2364;
32423: waveform_sig_loopback =-4112;
32424: waveform_sig_loopback =-6688;
32425: waveform_sig_loopback =-618;
32426: waveform_sig_loopback =-3287;
32427: waveform_sig_loopback =-4434;
32428: waveform_sig_loopback =-4352;
32429: waveform_sig_loopback =-3612;
32430: waveform_sig_loopback =-1488;
32431: waveform_sig_loopback =-3747;
32432: waveform_sig_loopback =-4895;
32433: waveform_sig_loopback =-2006;
32434: waveform_sig_loopback =-3920;
32435: waveform_sig_loopback =-2605;
32436: waveform_sig_loopback =-3576;
32437: waveform_sig_loopback =-3755;
32438: waveform_sig_loopback =-1570;
32439: waveform_sig_loopback =-4144;
32440: waveform_sig_loopback =-2885;
32441: waveform_sig_loopback =-2624;
32442: waveform_sig_loopback =-3052;
32443: waveform_sig_loopback =-3474;
32444: waveform_sig_loopback =-1925;
32445: waveform_sig_loopback =-2989;
32446: waveform_sig_loopback =-3618;
32447: waveform_sig_loopback =-1765;
32448: waveform_sig_loopback =-2786;
32449: waveform_sig_loopback =-3070;
32450: waveform_sig_loopback =-2684;
32451: waveform_sig_loopback =-1522;
32452: waveform_sig_loopback =-3329;
32453: waveform_sig_loopback =-3042;
32454: waveform_sig_loopback =-941;
32455: waveform_sig_loopback =-2771;
32456: waveform_sig_loopback =-3647;
32457: waveform_sig_loopback =-1127;
32458: waveform_sig_loopback =-1478;
32459: waveform_sig_loopback =-3720;
32460: waveform_sig_loopback =-2117;
32461: waveform_sig_loopback =-500;
32462: waveform_sig_loopback =-3490;
32463: waveform_sig_loopback =-409;
32464: waveform_sig_loopback =-2798;
32465: waveform_sig_loopback =-4573;
32466: waveform_sig_loopback =1149;
32467: waveform_sig_loopback =-1805;
32468: waveform_sig_loopback =-2384;
32469: waveform_sig_loopback =-2853;
32470: waveform_sig_loopback =-1668;
32471: waveform_sig_loopback =431;
32472: waveform_sig_loopback =-2456;
32473: waveform_sig_loopback =-2604;
32474: waveform_sig_loopback =-429;
32475: waveform_sig_loopback =-2221;
32476: waveform_sig_loopback =-365;
32477: waveform_sig_loopback =-2292;
32478: waveform_sig_loopback =-1574;
32479: waveform_sig_loopback =154;
32480: waveform_sig_loopback =-2673;
32481: waveform_sig_loopback =-540;
32482: waveform_sig_loopback =-1202;
32483: waveform_sig_loopback =-1128;
32484: waveform_sig_loopback =-1471;
32485: waveform_sig_loopback =-352;
32486: waveform_sig_loopback =-910;
32487: waveform_sig_loopback =-1880;
32488: waveform_sig_loopback =14;
32489: waveform_sig_loopback =-803;
32490: waveform_sig_loopback =-1381;
32491: waveform_sig_loopback =-658;
32492: waveform_sig_loopback =293;
32493: waveform_sig_loopback =-1569;
32494: waveform_sig_loopback =-1100;
32495: waveform_sig_loopback =980;
32496: waveform_sig_loopback =-1067;
32497: waveform_sig_loopback =-1791;
32498: waveform_sig_loopback =999;
32499: waveform_sig_loopback =73;
32500: waveform_sig_loopback =-1668;
32501: waveform_sig_loopback =-101;
32502: waveform_sig_loopback =1052;
32503: waveform_sig_loopback =-1258;
32504: waveform_sig_loopback =1304;
32505: waveform_sig_loopback =-1090;
32506: waveform_sig_loopback =-2182;
32507: waveform_sig_loopback =2594;
32508: waveform_sig_loopback =483;
32509: waveform_sig_loopback =-677;
32510: waveform_sig_loopback =-1159;
32511: waveform_sig_loopback =832;
32512: waveform_sig_loopback =1823;
32513: waveform_sig_loopback =-304;
32514: waveform_sig_loopback =-651;
32515: waveform_sig_loopback =1163;
32516: waveform_sig_loopback =143;
32517: waveform_sig_loopback =1211;
32518: waveform_sig_loopback =-455;
32519: waveform_sig_loopback =709;
32520: waveform_sig_loopback =1702;
32521: waveform_sig_loopback =-542;
32522: waveform_sig_loopback =1253;
32523: waveform_sig_loopback =639;
32524: waveform_sig_loopback =945;
32525: waveform_sig_loopback =305;
32526: waveform_sig_loopback =1637;
32527: waveform_sig_loopback =840;
32528: waveform_sig_loopback =146;
32529: waveform_sig_loopback =1830;
32530: waveform_sig_loopback =1179;
32531: waveform_sig_loopback =401;
32532: waveform_sig_loopback =1041;
32533: waveform_sig_loopback =2537;
32534: waveform_sig_loopback =-80;
32535: waveform_sig_loopback =1123;
32536: waveform_sig_loopback =2677;
32537: waveform_sig_loopback =528;
32538: waveform_sig_loopback =810;
32539: waveform_sig_loopback =2484;
32540: waveform_sig_loopback =1888;
32541: waveform_sig_loopback =388;
32542: waveform_sig_loopback =1629;
32543: waveform_sig_loopback =3204;
32544: waveform_sig_loopback =348;
32545: waveform_sig_loopback =3193;
32546: waveform_sig_loopback =949;
32547: waveform_sig_loopback =-634;
32548: waveform_sig_loopback =4686;
32549: waveform_sig_loopback =2314;
32550: waveform_sig_loopback =799;
32551: waveform_sig_loopback =1148;
32552: waveform_sig_loopback =2468;
32553: waveform_sig_loopback =3648;
32554: waveform_sig_loopback =1647;
32555: waveform_sig_loopback =991;
32556: waveform_sig_loopback =3191;
32557: waveform_sig_loopback =1931;
32558: waveform_sig_loopback =2945;
32559: waveform_sig_loopback =1484;
32560: waveform_sig_loopback =2570;
32561: waveform_sig_loopback =3367;
32562: waveform_sig_loopback =1434;
32563: waveform_sig_loopback =3032;
32564: waveform_sig_loopback =2352;
32565: waveform_sig_loopback =2895;
32566: waveform_sig_loopback =2002;
32567: waveform_sig_loopback =3423;
32568: waveform_sig_loopback =2766;
32569: waveform_sig_loopback =1736;
32570: waveform_sig_loopback =3842;
32571: waveform_sig_loopback =2983;
32572: waveform_sig_loopback =1935;
32573: waveform_sig_loopback =3533;
32574: waveform_sig_loopback =3758;
32575: waveform_sig_loopback =1706;
32576: waveform_sig_loopback =3334;
32577: waveform_sig_loopback =4185;
32578: waveform_sig_loopback =2530;
32579: waveform_sig_loopback =2306;
32580: waveform_sig_loopback =4269;
32581: waveform_sig_loopback =4023;
32582: waveform_sig_loopback =1713;
32583: waveform_sig_loopback =3549;
32584: waveform_sig_loopback =5097;
32585: waveform_sig_loopback =1796;
32586: waveform_sig_loopback =5353;
32587: waveform_sig_loopback =2209;
32588: waveform_sig_loopback =1332;
32589: waveform_sig_loopback =6818;
32590: waveform_sig_loopback =3502;
32591: waveform_sig_loopback =2721;
32592: waveform_sig_loopback =2930;
32593: waveform_sig_loopback =4161;
32594: waveform_sig_loopback =5415;
32595: waveform_sig_loopback =3088;
32596: waveform_sig_loopback =2864;
32597: waveform_sig_loopback =4943;
32598: waveform_sig_loopback =3592;
32599: waveform_sig_loopback =4459;
32600: waveform_sig_loopback =3299;
32601: waveform_sig_loopback =4347;
32602: waveform_sig_loopback =4820;
32603: waveform_sig_loopback =3330;
32604: waveform_sig_loopback =4448;
32605: waveform_sig_loopback =4222;
32606: waveform_sig_loopback =4628;
32607: waveform_sig_loopback =3171;
32608: waveform_sig_loopback =5675;
32609: waveform_sig_loopback =4041;
32610: waveform_sig_loopback =3416;
32611: waveform_sig_loopback =5768;
32612: waveform_sig_loopback =3944;
32613: waveform_sig_loopback =4118;
32614: waveform_sig_loopback =5014;
32615: waveform_sig_loopback =5080;
32616: waveform_sig_loopback =3637;
32617: waveform_sig_loopback =4656;
32618: waveform_sig_loopback =5982;
32619: waveform_sig_loopback =3851;
32620: waveform_sig_loopback =3862;
32621: waveform_sig_loopback =6067;
32622: waveform_sig_loopback =5331;
32623: waveform_sig_loopback =3234;
32624: waveform_sig_loopback =5264;
32625: waveform_sig_loopback =6665;
32626: waveform_sig_loopback =3075;
32627: waveform_sig_loopback =7128;
32628: waveform_sig_loopback =3469;
32629: waveform_sig_loopback =2901;
32630: waveform_sig_loopback =8544;
32631: waveform_sig_loopback =4506;
32632: waveform_sig_loopback =4398;
32633: waveform_sig_loopback =4543;
32634: waveform_sig_loopback =5295;
32635: waveform_sig_loopback =7196;
32636: waveform_sig_loopback =4274;
32637: waveform_sig_loopback =4376;
32638: waveform_sig_loopback =6578;
32639: waveform_sig_loopback =4586;
32640: waveform_sig_loopback =6184;
32641: waveform_sig_loopback =4670;
32642: waveform_sig_loopback =5504;
32643: waveform_sig_loopback =6470;
32644: waveform_sig_loopback =4564;
32645: waveform_sig_loopback =5788;
32646: waveform_sig_loopback =5781;
32647: waveform_sig_loopback =5576;
32648: waveform_sig_loopback =4875;
32649: waveform_sig_loopback =7022;
32650: waveform_sig_loopback =4927;
32651: waveform_sig_loopback =5206;
32652: waveform_sig_loopback =6899;
32653: waveform_sig_loopback =5254;
32654: waveform_sig_loopback =5504;
32655: waveform_sig_loopback =6131;
32656: waveform_sig_loopback =6479;
32657: waveform_sig_loopback =4974;
32658: waveform_sig_loopback =5819;
32659: waveform_sig_loopback =7256;
32660: waveform_sig_loopback =5109;
32661: waveform_sig_loopback =4997;
32662: waveform_sig_loopback =7497;
32663: waveform_sig_loopback =6352;
32664: waveform_sig_loopback =4355;
32665: waveform_sig_loopback =6859;
32666: waveform_sig_loopback =7333;
32667: waveform_sig_loopback =4462;
32668: waveform_sig_loopback =8559;
32669: waveform_sig_loopback =3906;
32670: waveform_sig_loopback =4768;
32671: waveform_sig_loopback =9504;
32672: waveform_sig_loopback =5416;
32673: waveform_sig_loopback =5940;
32674: waveform_sig_loopback =5154;
32675: waveform_sig_loopback =6850;
32676: waveform_sig_loopback =8330;
32677: waveform_sig_loopback =4822;
32678: waveform_sig_loopback =6048;
32679: waveform_sig_loopback =7321;
32680: waveform_sig_loopback =5644;
32681: waveform_sig_loopback =7535;
32682: waveform_sig_loopback =5265;
32683: waveform_sig_loopback =6911;
32684: waveform_sig_loopback =7406;
32685: waveform_sig_loopback =5300;
32686: waveform_sig_loopback =7163;
32687: waveform_sig_loopback =6569;
32688: waveform_sig_loopback =6496;
32689: waveform_sig_loopback =6084;
32690: waveform_sig_loopback =7794;
32691: waveform_sig_loopback =5880;
32692: waveform_sig_loopback =6334;
32693: waveform_sig_loopback =7575;
32694: waveform_sig_loopback =6261;
32695: waveform_sig_loopback =6500;
32696: waveform_sig_loopback =6845;
32697: waveform_sig_loopback =7540;
32698: waveform_sig_loopback =5702;
32699: waveform_sig_loopback =6635;
32700: waveform_sig_loopback =8423;
32701: waveform_sig_loopback =5533;
32702: waveform_sig_loopback =6047;
32703: waveform_sig_loopback =8536;
32704: waveform_sig_loopback =6644;
32705: waveform_sig_loopback =5575;
32706: waveform_sig_loopback =7583;
32707: waveform_sig_loopback =7803;
32708: waveform_sig_loopback =5749;
32709: waveform_sig_loopback =8871;
32710: waveform_sig_loopback =4644;
32711: waveform_sig_loopback =5932;
32712: waveform_sig_loopback =9699;
32713: waveform_sig_loopback =6555;
32714: waveform_sig_loopback =6338;
32715: waveform_sig_loopback =5723;
32716: waveform_sig_loopback =8017;
32717: waveform_sig_loopback =8480;
32718: waveform_sig_loopback =5676;
32719: waveform_sig_loopback =6827;
32720: waveform_sig_loopback =7621;
32721: waveform_sig_loopback =6648;
32722: waveform_sig_loopback =7961;
32723: waveform_sig_loopback =5736;
32724: waveform_sig_loopback =7831;
32725: waveform_sig_loopback =7710;
32726: waveform_sig_loopback =5972;
32727: waveform_sig_loopback =7819;
32728: waveform_sig_loopback =6944;
32729: waveform_sig_loopback =7075;
32730: waveform_sig_loopback =6781;
32731: waveform_sig_loopback =8030;
32732: waveform_sig_loopback =6486;
32733: waveform_sig_loopback =6901;
32734: waveform_sig_loopback =7739;
32735: waveform_sig_loopback =7176;
32736: waveform_sig_loopback =6460;
32737: waveform_sig_loopback =7487;
32738: waveform_sig_loopback =8146;
32739: waveform_sig_loopback =5521;
32740: waveform_sig_loopback =7659;
32741: waveform_sig_loopback =8492;
32742: waveform_sig_loopback =5773;
32743: waveform_sig_loopback =6885;
32744: waveform_sig_loopback =8454;
32745: waveform_sig_loopback =7140;
32746: waveform_sig_loopback =5947;
32747: waveform_sig_loopback =7716;
32748: waveform_sig_loopback =8307;
32749: waveform_sig_loopback =5949;
32750: waveform_sig_loopback =9098;
32751: waveform_sig_loopback =5006;
32752: waveform_sig_loopback =6197;
32753: waveform_sig_loopback =9986;
32754: waveform_sig_loopback =6910;
32755: waveform_sig_loopback =6226;
32756: waveform_sig_loopback =6266;
32757: waveform_sig_loopback =8264;
32758: waveform_sig_loopback =8403;
32759: waveform_sig_loopback =6092;
32760: waveform_sig_loopback =6865;
32761: waveform_sig_loopback =7754;
32762: waveform_sig_loopback =7004;
32763: waveform_sig_loopback =7787;
32764: waveform_sig_loopback =6028;
32765: waveform_sig_loopback =8097;
32766: waveform_sig_loopback =7415;
32767: waveform_sig_loopback =6372;

default: waveform_sig_loopback= 0;
endcase

case(msg_count_tx_idx)
0: waveform_sig_rx =-319;
1: waveform_sig_rx =-702;
2: waveform_sig_rx =-689;
3: waveform_sig_rx =-376;
4: waveform_sig_rx =-605;
5: waveform_sig_rx =-701;
6: waveform_sig_rx =-447;
7: waveform_sig_rx =-501;
8: waveform_sig_rx =-584;
9: waveform_sig_rx =-608;
10: waveform_sig_rx =-364;
11: waveform_sig_rx =-565;
12: waveform_sig_rx =-665;
13: waveform_sig_rx =-311;
14: waveform_sig_rx =-543;
15: waveform_sig_rx =-628;
16: waveform_sig_rx =-388;
17: waveform_sig_rx =-393;
18: waveform_sig_rx =-663;
19: waveform_sig_rx =-434;
20: waveform_sig_rx =-314;
21: waveform_sig_rx =-627;
22: waveform_sig_rx =-459;
23: waveform_sig_rx =-325;
24: waveform_sig_rx =-525;
25: waveform_sig_rx =-441;
26: waveform_sig_rx =-451;
27: waveform_sig_rx =-425;
28: waveform_sig_rx =-374;
29: waveform_sig_rx =-484;
30: waveform_sig_rx =-288;
31: waveform_sig_rx =-606;
32: waveform_sig_rx =-164;
33: waveform_sig_rx =-464;
34: waveform_sig_rx =-492;
35: waveform_sig_rx =-120;
36: waveform_sig_rx =-535;
37: waveform_sig_rx =-420;
38: waveform_sig_rx =-85;
39: waveform_sig_rx =-513;
40: waveform_sig_rx =-397;
41: waveform_sig_rx =-75;
42: waveform_sig_rx =-465;
43: waveform_sig_rx =-337;
44: waveform_sig_rx =-165;
45: waveform_sig_rx =-283;
46: waveform_sig_rx =-421;
47: waveform_sig_rx =-195;
48: waveform_sig_rx =-193;
49: waveform_sig_rx =-377;
50: waveform_sig_rx =-301;
51: waveform_sig_rx =-79;
52: waveform_sig_rx =-329;
53: waveform_sig_rx =-359;
54: waveform_sig_rx =-31;
55: waveform_sig_rx =-263;
56: waveform_sig_rx =-348;
57: waveform_sig_rx =-53;
58: waveform_sig_rx =-143;
59: waveform_sig_rx =-342;
60: waveform_sig_rx =-120;
61: waveform_sig_rx =-112;
62: waveform_sig_rx =-283;
63: waveform_sig_rx =-194;
64: waveform_sig_rx =-25;
65: waveform_sig_rx =-194;
66: waveform_sig_rx =-208;
67: waveform_sig_rx =-88;
68: waveform_sig_rx =-155;
69: waveform_sig_rx =-128;
70: waveform_sig_rx =-113;
71: waveform_sig_rx =-56;
72: waveform_sig_rx =-293;
73: waveform_sig_rx =158;
74: waveform_sig_rx =-275;
75: waveform_sig_rx =-131;
76: waveform_sig_rx =163;
77: waveform_sig_rx =-279;
78: waveform_sig_rx =-53;
79: waveform_sig_rx =170;
80: waveform_sig_rx =-197;
81: waveform_sig_rx =-77;
82: waveform_sig_rx =177;
83: waveform_sig_rx =-152;
84: waveform_sig_rx =-72;
85: waveform_sig_rx =99;
86: waveform_sig_rx =2;
87: waveform_sig_rx =-172;
88: waveform_sig_rx =89;
89: waveform_sig_rx =102;
90: waveform_sig_rx =-104;
91: waveform_sig_rx =-8;
92: waveform_sig_rx =236;
93: waveform_sig_rx =-87;
94: waveform_sig_rx =-34;
95: waveform_sig_rx =270;
96: waveform_sig_rx =-29;
97: waveform_sig_rx =-5;
98: waveform_sig_rx =202;
99: waveform_sig_rx =120;
100: waveform_sig_rx =-31;
101: waveform_sig_rx =115;
102: waveform_sig_rx =231;
103: waveform_sig_rx =-1;
104: waveform_sig_rx =59;
105: waveform_sig_rx =351;
106: waveform_sig_rx =18;
107: waveform_sig_rx =110;
108: waveform_sig_rx =225;
109: waveform_sig_rx =97;
110: waveform_sig_rx =210;
111: waveform_sig_rx =168;
112: waveform_sig_rx =195;
113: waveform_sig_rx =54;
114: waveform_sig_rx =417;
115: waveform_sig_rx =10;
116: waveform_sig_rx =198;
117: waveform_sig_rx =403;
118: waveform_sig_rx =17;
119: waveform_sig_rx =254;
120: waveform_sig_rx =415;
121: waveform_sig_rx =79;
122: waveform_sig_rx =220;
123: waveform_sig_rx =436;
124: waveform_sig_rx =157;
125: waveform_sig_rx =229;
126: waveform_sig_rx =382;
127: waveform_sig_rx =330;
128: waveform_sig_rx =93;
129: waveform_sig_rx =442;
130: waveform_sig_rx =384;
131: waveform_sig_rx =157;
132: waveform_sig_rx =352;
133: waveform_sig_rx =479;
134: waveform_sig_rx =205;
135: waveform_sig_rx =310;
136: waveform_sig_rx =478;
137: waveform_sig_rx =301;
138: waveform_sig_rx =266;
139: waveform_sig_rx =461;
140: waveform_sig_rx =469;
141: waveform_sig_rx =215;
142: waveform_sig_rx =445;
143: waveform_sig_rx =534;
144: waveform_sig_rx =233;
145: waveform_sig_rx =378;
146: waveform_sig_rx =623;
147: waveform_sig_rx =276;
148: waveform_sig_rx =445;
149: waveform_sig_rx =481;
150: waveform_sig_rx =364;
151: waveform_sig_rx =528;
152: waveform_sig_rx =421;
153: waveform_sig_rx =478;
154: waveform_sig_rx =356;
155: waveform_sig_rx =675;
156: waveform_sig_rx =297;
157: waveform_sig_rx =499;
158: waveform_sig_rx =645;
159: waveform_sig_rx =324;
160: waveform_sig_rx =527;
161: waveform_sig_rx =671;
162: waveform_sig_rx =376;
163: waveform_sig_rx =463;
164: waveform_sig_rx =730;
165: waveform_sig_rx =435;
166: waveform_sig_rx =468;
167: waveform_sig_rx =709;
168: waveform_sig_rx =570;
169: waveform_sig_rx =334;
170: waveform_sig_rx =752;
171: waveform_sig_rx =600;
172: waveform_sig_rx =458;
173: waveform_sig_rx =643;
174: waveform_sig_rx =706;
175: waveform_sig_rx =511;
176: waveform_sig_rx =550;
177: waveform_sig_rx =747;
178: waveform_sig_rx =592;
179: waveform_sig_rx =493;
180: waveform_sig_rx =771;
181: waveform_sig_rx =709;
182: waveform_sig_rx =458;
183: waveform_sig_rx =749;
184: waveform_sig_rx =764;
185: waveform_sig_rx =486;
186: waveform_sig_rx =655;
187: waveform_sig_rx =861;
188: waveform_sig_rx =509;
189: waveform_sig_rx =727;
190: waveform_sig_rx =685;
191: waveform_sig_rx =631;
192: waveform_sig_rx =791;
193: waveform_sig_rx =648;
194: waveform_sig_rx =747;
195: waveform_sig_rx =603;
196: waveform_sig_rx =891;
197: waveform_sig_rx =596;
198: waveform_sig_rx =710;
199: waveform_sig_rx =922;
200: waveform_sig_rx =591;
201: waveform_sig_rx =720;
202: waveform_sig_rx =993;
203: waveform_sig_rx =577;
204: waveform_sig_rx =739;
205: waveform_sig_rx =1008;
206: waveform_sig_rx =603;
207: waveform_sig_rx =779;
208: waveform_sig_rx =919;
209: waveform_sig_rx =782;
210: waveform_sig_rx =620;
211: waveform_sig_rx =968;
212: waveform_sig_rx =818;
213: waveform_sig_rx =700;
214: waveform_sig_rx =859;
215: waveform_sig_rx =922;
216: waveform_sig_rx =756;
217: waveform_sig_rx =782;
218: waveform_sig_rx =976;
219: waveform_sig_rx =833;
220: waveform_sig_rx =678;
221: waveform_sig_rx =1032;
222: waveform_sig_rx =890;
223: waveform_sig_rx =646;
224: waveform_sig_rx =1036;
225: waveform_sig_rx =929;
226: waveform_sig_rx =740;
227: waveform_sig_rx =929;
228: waveform_sig_rx =1021;
229: waveform_sig_rx =769;
230: waveform_sig_rx =918;
231: waveform_sig_rx =867;
232: waveform_sig_rx =915;
233: waveform_sig_rx =935;
234: waveform_sig_rx =874;
235: waveform_sig_rx =975;
236: waveform_sig_rx =770;
237: waveform_sig_rx =1142;
238: waveform_sig_rx =770;
239: waveform_sig_rx =904;
240: waveform_sig_rx =1140;
241: waveform_sig_rx =728;
242: waveform_sig_rx =969;
243: waveform_sig_rx =1185;
244: waveform_sig_rx =722;
245: waveform_sig_rx =967;
246: waveform_sig_rx =1192;
247: waveform_sig_rx =768;
248: waveform_sig_rx =983;
249: waveform_sig_rx =1103;
250: waveform_sig_rx =932;
251: waveform_sig_rx =831;
252: waveform_sig_rx =1146;
253: waveform_sig_rx =973;
254: waveform_sig_rx =896;
255: waveform_sig_rx =990;
256: waveform_sig_rx =1126;
257: waveform_sig_rx =901;
258: waveform_sig_rx =914;
259: waveform_sig_rx =1202;
260: waveform_sig_rx =924;
261: waveform_sig_rx =872;
262: waveform_sig_rx =1234;
263: waveform_sig_rx =977;
264: waveform_sig_rx =867;
265: waveform_sig_rx =1179;
266: waveform_sig_rx =1048;
267: waveform_sig_rx =935;
268: waveform_sig_rx =1043;
269: waveform_sig_rx =1184;
270: waveform_sig_rx =923;
271: waveform_sig_rx =1032;
272: waveform_sig_rx =1058;
273: waveform_sig_rx =1044;
274: waveform_sig_rx =1066;
275: waveform_sig_rx =1073;
276: waveform_sig_rx =1071;
277: waveform_sig_rx =946;
278: waveform_sig_rx =1297;
279: waveform_sig_rx =844;
280: waveform_sig_rx =1095;
281: waveform_sig_rx =1269;
282: waveform_sig_rx =843;
283: waveform_sig_rx =1140;
284: waveform_sig_rx =1288;
285: waveform_sig_rx =841;
286: waveform_sig_rx =1146;
287: waveform_sig_rx =1275;
288: waveform_sig_rx =872;
289: waveform_sig_rx =1127;
290: waveform_sig_rx =1187;
291: waveform_sig_rx =1065;
292: waveform_sig_rx =965;
293: waveform_sig_rx =1236;
294: waveform_sig_rx =1125;
295: waveform_sig_rx =1007;
296: waveform_sig_rx =1124;
297: waveform_sig_rx =1294;
298: waveform_sig_rx =938;
299: waveform_sig_rx =1094;
300: waveform_sig_rx =1296;
301: waveform_sig_rx =972;
302: waveform_sig_rx =1066;
303: waveform_sig_rx =1263;
304: waveform_sig_rx =1095;
305: waveform_sig_rx =989;
306: waveform_sig_rx =1219;
307: waveform_sig_rx =1183;
308: waveform_sig_rx =991;
309: waveform_sig_rx =1138;
310: waveform_sig_rx =1307;
311: waveform_sig_rx =975;
312: waveform_sig_rx =1172;
313: waveform_sig_rx =1134;
314: waveform_sig_rx =1136;
315: waveform_sig_rx =1141;
316: waveform_sig_rx =1175;
317: waveform_sig_rx =1091;
318: waveform_sig_rx =1050;
319: waveform_sig_rx =1376;
320: waveform_sig_rx =902;
321: waveform_sig_rx =1227;
322: waveform_sig_rx =1269;
323: waveform_sig_rx =896;
324: waveform_sig_rx =1265;
325: waveform_sig_rx =1266;
326: waveform_sig_rx =934;
327: waveform_sig_rx =1203;
328: waveform_sig_rx =1281;
329: waveform_sig_rx =990;
330: waveform_sig_rx =1141;
331: waveform_sig_rx =1262;
332: waveform_sig_rx =1122;
333: waveform_sig_rx =992;
334: waveform_sig_rx =1324;
335: waveform_sig_rx =1154;
336: waveform_sig_rx =1003;
337: waveform_sig_rx =1188;
338: waveform_sig_rx =1273;
339: waveform_sig_rx =957;
340: waveform_sig_rx =1174;
341: waveform_sig_rx =1283;
342: waveform_sig_rx =1013;
343: waveform_sig_rx =1110;
344: waveform_sig_rx =1266;
345: waveform_sig_rx =1140;
346: waveform_sig_rx =1022;
347: waveform_sig_rx =1220;
348: waveform_sig_rx =1250;
349: waveform_sig_rx =976;
350: waveform_sig_rx =1172;
351: waveform_sig_rx =1338;
352: waveform_sig_rx =940;
353: waveform_sig_rx =1238;
354: waveform_sig_rx =1110;
355: waveform_sig_rx =1126;
356: waveform_sig_rx =1190;
357: waveform_sig_rx =1162;
358: waveform_sig_rx =1088;
359: waveform_sig_rx =1094;
360: waveform_sig_rx =1324;
361: waveform_sig_rx =904;
362: waveform_sig_rx =1255;
363: waveform_sig_rx =1212;
364: waveform_sig_rx =923;
365: waveform_sig_rx =1250;
366: waveform_sig_rx =1220;
367: waveform_sig_rx =949;
368: waveform_sig_rx =1167;
369: waveform_sig_rx =1262;
370: waveform_sig_rx =984;
371: waveform_sig_rx =1099;
372: waveform_sig_rx =1254;
373: waveform_sig_rx =1061;
374: waveform_sig_rx =947;
375: waveform_sig_rx =1321;
376: waveform_sig_rx =1061;
377: waveform_sig_rx =998;
378: waveform_sig_rx =1197;
379: waveform_sig_rx =1208;
380: waveform_sig_rx =969;
381: waveform_sig_rx =1171;
382: waveform_sig_rx =1206;
383: waveform_sig_rx =1003;
384: waveform_sig_rx =1023;
385: waveform_sig_rx =1203;
386: waveform_sig_rx =1109;
387: waveform_sig_rx =904;
388: waveform_sig_rx =1230;
389: waveform_sig_rx =1165;
390: waveform_sig_rx =885;
391: waveform_sig_rx =1171;
392: waveform_sig_rx =1204;
393: waveform_sig_rx =895;
394: waveform_sig_rx =1196;
395: waveform_sig_rx =980;
396: waveform_sig_rx =1110;
397: waveform_sig_rx =1065;
398: waveform_sig_rx =1074;
399: waveform_sig_rx =1029;
400: waveform_sig_rx =1034;
401: waveform_sig_rx =1241;
402: waveform_sig_rx =842;
403: waveform_sig_rx =1177;
404: waveform_sig_rx =1128;
405: waveform_sig_rx =876;
406: waveform_sig_rx =1151;
407: waveform_sig_rx =1157;
408: waveform_sig_rx =887;
409: waveform_sig_rx =1035;
410: waveform_sig_rx =1219;
411: waveform_sig_rx =842;
412: waveform_sig_rx =1020;
413: waveform_sig_rx =1226;
414: waveform_sig_rx =882;
415: waveform_sig_rx =919;
416: waveform_sig_rx =1222;
417: waveform_sig_rx =897;
418: waveform_sig_rx =973;
419: waveform_sig_rx =1033;
420: waveform_sig_rx =1101;
421: waveform_sig_rx =871;
422: waveform_sig_rx =980;
423: waveform_sig_rx =1133;
424: waveform_sig_rx =870;
425: waveform_sig_rx =900;
426: waveform_sig_rx =1137;
427: waveform_sig_rx =941;
428: waveform_sig_rx =801;
429: waveform_sig_rx =1121;
430: waveform_sig_rx =980;
431: waveform_sig_rx =805;
432: waveform_sig_rx =1072;
433: waveform_sig_rx =1038;
434: waveform_sig_rx =792;
435: waveform_sig_rx =1053;
436: waveform_sig_rx =837;
437: waveform_sig_rx =980;
438: waveform_sig_rx =905;
439: waveform_sig_rx =957;
440: waveform_sig_rx =869;
441: waveform_sig_rx =879;
442: waveform_sig_rx =1054;
443: waveform_sig_rx =701;
444: waveform_sig_rx =993;
445: waveform_sig_rx =990;
446: waveform_sig_rx =716;
447: waveform_sig_rx =961;
448: waveform_sig_rx =1049;
449: waveform_sig_rx =622;
450: waveform_sig_rx =911;
451: waveform_sig_rx =1072;
452: waveform_sig_rx =607;
453: waveform_sig_rx =947;
454: waveform_sig_rx =995;
455: waveform_sig_rx =700;
456: waveform_sig_rx =818;
457: waveform_sig_rx =971;
458: waveform_sig_rx =784;
459: waveform_sig_rx =780;
460: waveform_sig_rx =814;
461: waveform_sig_rx =981;
462: waveform_sig_rx =622;
463: waveform_sig_rx =843;
464: waveform_sig_rx =951;
465: waveform_sig_rx =639;
466: waveform_sig_rx =757;
467: waveform_sig_rx =922;
468: waveform_sig_rx =753;
469: waveform_sig_rx =615;
470: waveform_sig_rx =953;
471: waveform_sig_rx =781;
472: waveform_sig_rx =588;
473: waveform_sig_rx =903;
474: waveform_sig_rx =789;
475: waveform_sig_rx =631;
476: waveform_sig_rx =831;
477: waveform_sig_rx =602;
478: waveform_sig_rx =878;
479: waveform_sig_rx =631;
480: waveform_sig_rx =799;
481: waveform_sig_rx =682;
482: waveform_sig_rx =634;
483: waveform_sig_rx =910;
484: waveform_sig_rx =453;
485: waveform_sig_rx =791;
486: waveform_sig_rx =803;
487: waveform_sig_rx =408;
488: waveform_sig_rx =833;
489: waveform_sig_rx =747;
490: waveform_sig_rx =411;
491: waveform_sig_rx =762;
492: waveform_sig_rx =746;
493: waveform_sig_rx =430;
494: waveform_sig_rx =700;
495: waveform_sig_rx =758;
496: waveform_sig_rx =497;
497: waveform_sig_rx =546;
498: waveform_sig_rx =763;
499: waveform_sig_rx =546;
500: waveform_sig_rx =548;
501: waveform_sig_rx =608;
502: waveform_sig_rx =728;
503: waveform_sig_rx =385;
504: waveform_sig_rx =630;
505: waveform_sig_rx =731;
506: waveform_sig_rx =383;
507: waveform_sig_rx =545;
508: waveform_sig_rx =722;
509: waveform_sig_rx =444;
510: waveform_sig_rx =448;
511: waveform_sig_rx =701;
512: waveform_sig_rx =481;
513: waveform_sig_rx =418;
514: waveform_sig_rx =575;
515: waveform_sig_rx =585;
516: waveform_sig_rx =399;
517: waveform_sig_rx =521;
518: waveform_sig_rx =432;
519: waveform_sig_rx =550;
520: waveform_sig_rx =371;
521: waveform_sig_rx =594;
522: waveform_sig_rx =302;
523: waveform_sig_rx =436;
524: waveform_sig_rx =650;
525: waveform_sig_rx =122;
526: waveform_sig_rx =630;
527: waveform_sig_rx =456;
528: waveform_sig_rx =191;
529: waveform_sig_rx =595;
530: waveform_sig_rx =439;
531: waveform_sig_rx =211;
532: waveform_sig_rx =498;
533: waveform_sig_rx =489;
534: waveform_sig_rx =177;
535: waveform_sig_rx =460;
536: waveform_sig_rx =459;
537: waveform_sig_rx =231;
538: waveform_sig_rx =309;
539: waveform_sig_rx =456;
540: waveform_sig_rx =301;
541: waveform_sig_rx =234;
542: waveform_sig_rx =364;
543: waveform_sig_rx =482;
544: waveform_sig_rx =48;
545: waveform_sig_rx =408;
546: waveform_sig_rx =425;
547: waveform_sig_rx =75;
548: waveform_sig_rx =335;
549: waveform_sig_rx =365;
550: waveform_sig_rx =175;
551: waveform_sig_rx =187;
552: waveform_sig_rx =332;
553: waveform_sig_rx =270;
554: waveform_sig_rx =84;
555: waveform_sig_rx =307;
556: waveform_sig_rx =364;
557: waveform_sig_rx =-4;
558: waveform_sig_rx =305;
559: waveform_sig_rx =140;
560: waveform_sig_rx =216;
561: waveform_sig_rx =164;
562: waveform_sig_rx =258;
563: waveform_sig_rx =4;
564: waveform_sig_rx =229;
565: waveform_sig_rx =258;
566: waveform_sig_rx =-115;
567: waveform_sig_rx =329;
568: waveform_sig_rx =121;
569: waveform_sig_rx =-79;
570: waveform_sig_rx =307;
571: waveform_sig_rx =134;
572: waveform_sig_rx =-105;
573: waveform_sig_rx =233;
574: waveform_sig_rx =132;
575: waveform_sig_rx =-93;
576: waveform_sig_rx =130;
577: waveform_sig_rx =125;
578: waveform_sig_rx =-17;
579: waveform_sig_rx =-78;
580: waveform_sig_rx =218;
581: waveform_sig_rx =-34;
582: waveform_sig_rx =-122;
583: waveform_sig_rx =154;
584: waveform_sig_rx =49;
585: waveform_sig_rx =-227;
586: waveform_sig_rx =132;
587: waveform_sig_rx =6;
588: waveform_sig_rx =-133;
589: waveform_sig_rx =-47;
590: waveform_sig_rx =92;
591: waveform_sig_rx =-74;
592: waveform_sig_rx =-190;
593: waveform_sig_rx =96;
594: waveform_sig_rx =-55;
595: waveform_sig_rx =-268;
596: waveform_sig_rx =38;
597: waveform_sig_rx =-4;
598: waveform_sig_rx =-296;
599: waveform_sig_rx =23;
600: waveform_sig_rx =-196;
601: waveform_sig_rx =-74;
602: waveform_sig_rx =-127;
603: waveform_sig_rx =-89;
604: waveform_sig_rx =-273;
605: waveform_sig_rx =-73;
606: waveform_sig_rx =-86;
607: waveform_sig_rx =-384;
608: waveform_sig_rx =13;
609: waveform_sig_rx =-217;
610: waveform_sig_rx =-334;
611: waveform_sig_rx =-37;
612: waveform_sig_rx =-184;
613: waveform_sig_rx =-399;
614: waveform_sig_rx =-115;
615: waveform_sig_rx =-154;
616: waveform_sig_rx =-410;
617: waveform_sig_rx =-200;
618: waveform_sig_rx =-109;
619: waveform_sig_rx =-397;
620: waveform_sig_rx =-358;
621: waveform_sig_rx =-38;
622: waveform_sig_rx =-409;
623: waveform_sig_rx =-352;
624: waveform_sig_rx =-188;
625: waveform_sig_rx =-284;
626: waveform_sig_rx =-460;
627: waveform_sig_rx =-234;
628: waveform_sig_rx =-262;
629: waveform_sig_rx =-429;
630: waveform_sig_rx =-381;
631: waveform_sig_rx =-164;
632: waveform_sig_rx =-426;
633: waveform_sig_rx =-500;
634: waveform_sig_rx =-160;
635: waveform_sig_rx =-411;
636: waveform_sig_rx =-551;
637: waveform_sig_rx =-228;
638: waveform_sig_rx =-341;
639: waveform_sig_rx =-568;
640: waveform_sig_rx =-258;
641: waveform_sig_rx =-551;
642: waveform_sig_rx =-339;
643: waveform_sig_rx =-459;
644: waveform_sig_rx =-394;
645: waveform_sig_rx =-537;
646: waveform_sig_rx =-400;
647: waveform_sig_rx =-387;
648: waveform_sig_rx =-644;
649: waveform_sig_rx =-322;
650: waveform_sig_rx =-472;
651: waveform_sig_rx =-636;
652: waveform_sig_rx =-371;
653: waveform_sig_rx =-412;
654: waveform_sig_rx =-738;
655: waveform_sig_rx =-381;
656: waveform_sig_rx =-425;
657: waveform_sig_rx =-760;
658: waveform_sig_rx =-434;
659: waveform_sig_rx =-413;
660: waveform_sig_rx =-725;
661: waveform_sig_rx =-577;
662: waveform_sig_rx =-392;
663: waveform_sig_rx =-691;
664: waveform_sig_rx =-601;
665: waveform_sig_rx =-513;
666: waveform_sig_rx =-537;
667: waveform_sig_rx =-736;
668: waveform_sig_rx =-547;
669: waveform_sig_rx =-485;
670: waveform_sig_rx =-732;
671: waveform_sig_rx =-650;
672: waveform_sig_rx =-395;
673: waveform_sig_rx =-759;
674: waveform_sig_rx =-734;
675: waveform_sig_rx =-422;
676: waveform_sig_rx =-734;
677: waveform_sig_rx =-753;
678: waveform_sig_rx =-509;
679: waveform_sig_rx =-647;
680: waveform_sig_rx =-781;
681: waveform_sig_rx =-575;
682: waveform_sig_rx =-800;
683: waveform_sig_rx =-570;
684: waveform_sig_rx =-782;
685: waveform_sig_rx =-622;
686: waveform_sig_rx =-798;
687: waveform_sig_rx =-659;
688: waveform_sig_rx =-628;
689: waveform_sig_rx =-926;
690: waveform_sig_rx =-591;
691: waveform_sig_rx =-701;
692: waveform_sig_rx =-964;
693: waveform_sig_rx =-567;
694: waveform_sig_rx =-702;
695: waveform_sig_rx =-1043;
696: waveform_sig_rx =-556;
697: waveform_sig_rx =-723;
698: waveform_sig_rx =-991;
699: waveform_sig_rx =-663;
700: waveform_sig_rx =-719;
701: waveform_sig_rx =-967;
702: waveform_sig_rx =-796;
703: waveform_sig_rx =-673;
704: waveform_sig_rx =-898;
705: waveform_sig_rx =-859;
706: waveform_sig_rx =-778;
707: waveform_sig_rx =-733;
708: waveform_sig_rx =-1018;
709: waveform_sig_rx =-763;
710: waveform_sig_rx =-719;
711: waveform_sig_rx =-1048;
712: waveform_sig_rx =-831;
713: waveform_sig_rx =-677;
714: waveform_sig_rx =-1049;
715: waveform_sig_rx =-889;
716: waveform_sig_rx =-718;
717: waveform_sig_rx =-977;
718: waveform_sig_rx =-966;
719: waveform_sig_rx =-782;
720: waveform_sig_rx =-831;
721: waveform_sig_rx =-1022;
722: waveform_sig_rx =-826;
723: waveform_sig_rx =-1001;
724: waveform_sig_rx =-830;
725: waveform_sig_rx =-1008;
726: waveform_sig_rx =-827;
727: waveform_sig_rx =-1079;
728: waveform_sig_rx =-861;
729: waveform_sig_rx =-841;
730: waveform_sig_rx =-1166;
731: waveform_sig_rx =-758;
732: waveform_sig_rx =-912;
733: waveform_sig_rx =-1198;
734: waveform_sig_rx =-707;
735: waveform_sig_rx =-969;
736: waveform_sig_rx =-1227;
737: waveform_sig_rx =-711;
738: waveform_sig_rx =-1021;
739: waveform_sig_rx =-1137;
740: waveform_sig_rx =-857;
741: waveform_sig_rx =-966;
742: waveform_sig_rx =-1089;
743: waveform_sig_rx =-1029;
744: waveform_sig_rx =-858;
745: waveform_sig_rx =-1062;
746: waveform_sig_rx =-1110;
747: waveform_sig_rx =-907;
748: waveform_sig_rx =-951;
749: waveform_sig_rx =-1233;
750: waveform_sig_rx =-888;
751: waveform_sig_rx =-945;
752: waveform_sig_rx =-1235;
753: waveform_sig_rx =-979;
754: waveform_sig_rx =-887;
755: waveform_sig_rx =-1214;
756: waveform_sig_rx =-1055;
757: waveform_sig_rx =-943;
758: waveform_sig_rx =-1108;
759: waveform_sig_rx =-1139;
760: waveform_sig_rx =-972;
761: waveform_sig_rx =-976;
762: waveform_sig_rx =-1217;
763: waveform_sig_rx =-977;
764: waveform_sig_rx =-1119;
765: waveform_sig_rx =-1025;
766: waveform_sig_rx =-1126;
767: waveform_sig_rx =-972;
768: waveform_sig_rx =-1267;
769: waveform_sig_rx =-945;
770: waveform_sig_rx =-1046;
771: waveform_sig_rx =-1310;
772: waveform_sig_rx =-839;
773: waveform_sig_rx =-1155;
774: waveform_sig_rx =-1279;
775: waveform_sig_rx =-840;
776: waveform_sig_rx =-1172;
777: waveform_sig_rx =-1271;
778: waveform_sig_rx =-873;
779: waveform_sig_rx =-1159;
780: waveform_sig_rx =-1203;
781: waveform_sig_rx =-1029;
782: waveform_sig_rx =-1044;
783: waveform_sig_rx =-1218;
784: waveform_sig_rx =-1155;
785: waveform_sig_rx =-948;
786: waveform_sig_rx =-1210;
787: waveform_sig_rx =-1229;
788: waveform_sig_rx =-974;
789: waveform_sig_rx =-1103;
790: waveform_sig_rx =-1325;
791: waveform_sig_rx =-965;
792: waveform_sig_rx =-1106;
793: waveform_sig_rx =-1305;
794: waveform_sig_rx =-1064;
795: waveform_sig_rx =-1031;
796: waveform_sig_rx =-1264;
797: waveform_sig_rx =-1168;
798: waveform_sig_rx =-1022;
799: waveform_sig_rx =-1165;
800: waveform_sig_rx =-1283;
801: waveform_sig_rx =-993;
802: waveform_sig_rx =-1084;
803: waveform_sig_rx =-1329;
804: waveform_sig_rx =-985;
805: waveform_sig_rx =-1245;
806: waveform_sig_rx =-1109;
807: waveform_sig_rx =-1146;
808: waveform_sig_rx =-1088;
809: waveform_sig_rx =-1318;
810: waveform_sig_rx =-985;
811: waveform_sig_rx =-1196;
812: waveform_sig_rx =-1304;
813: waveform_sig_rx =-924;
814: waveform_sig_rx =-1253;
815: waveform_sig_rx =-1252;
816: waveform_sig_rx =-946;
817: waveform_sig_rx =-1210;
818: waveform_sig_rx =-1314;
819: waveform_sig_rx =-975;
820: waveform_sig_rx =-1186;
821: waveform_sig_rx =-1272;
822: waveform_sig_rx =-1075;
823: waveform_sig_rx =-1064;
824: waveform_sig_rx =-1308;
825: waveform_sig_rx =-1191;
826: waveform_sig_rx =-980;
827: waveform_sig_rx =-1296;
828: waveform_sig_rx =-1234;
829: waveform_sig_rx =-991;
830: waveform_sig_rx =-1197;
831: waveform_sig_rx =-1299;
832: waveform_sig_rx =-991;
833: waveform_sig_rx =-1176;
834: waveform_sig_rx =-1250;
835: waveform_sig_rx =-1125;
836: waveform_sig_rx =-1039;
837: waveform_sig_rx =-1249;
838: waveform_sig_rx =-1248;
839: waveform_sig_rx =-947;
840: waveform_sig_rx =-1222;
841: waveform_sig_rx =-1303;
842: waveform_sig_rx =-934;
843: waveform_sig_rx =-1190;
844: waveform_sig_rx =-1260;
845: waveform_sig_rx =-1015;
846: waveform_sig_rx =-1297;
847: waveform_sig_rx =-1041;
848: waveform_sig_rx =-1199;
849: waveform_sig_rx =-1077;
850: waveform_sig_rx =-1281;
851: waveform_sig_rx =-975;
852: waveform_sig_rx =-1169;
853: waveform_sig_rx =-1257;
854: waveform_sig_rx =-925;
855: waveform_sig_rx =-1222;
856: waveform_sig_rx =-1207;
857: waveform_sig_rx =-948;
858: waveform_sig_rx =-1166;
859: waveform_sig_rx =-1259;
860: waveform_sig_rx =-957;
861: waveform_sig_rx =-1097;
862: waveform_sig_rx =-1272;
863: waveform_sig_rx =-1027;
864: waveform_sig_rx =-1005;
865: waveform_sig_rx =-1338;
866: waveform_sig_rx =-1038;
867: waveform_sig_rx =-957;
868: waveform_sig_rx =-1262;
869: waveform_sig_rx =-1099;
870: waveform_sig_rx =-996;
871: waveform_sig_rx =-1123;
872: waveform_sig_rx =-1224;
873: waveform_sig_rx =-970;
874: waveform_sig_rx =-1056;
875: waveform_sig_rx =-1216;
876: waveform_sig_rx =-1056;
877: waveform_sig_rx =-932;
878: waveform_sig_rx =-1225;
879: waveform_sig_rx =-1136;
880: waveform_sig_rx =-879;
881: waveform_sig_rx =-1217;
882: waveform_sig_rx =-1182;
883: waveform_sig_rx =-870;
884: waveform_sig_rx =-1153;
885: waveform_sig_rx =-1118;
886: waveform_sig_rx =-969;
887: waveform_sig_rx =-1190;
888: waveform_sig_rx =-922;
889: waveform_sig_rx =-1139;
890: waveform_sig_rx =-949;
891: waveform_sig_rx =-1197;
892: waveform_sig_rx =-896;
893: waveform_sig_rx =-1056;
894: waveform_sig_rx =-1163;
895: waveform_sig_rx =-850;
896: waveform_sig_rx =-1093;
897: waveform_sig_rx =-1130;
898: waveform_sig_rx =-829;
899: waveform_sig_rx =-1033;
900: waveform_sig_rx =-1203;
901: waveform_sig_rx =-791;
902: waveform_sig_rx =-1029;
903: waveform_sig_rx =-1185;
904: waveform_sig_rx =-802;
905: waveform_sig_rx =-953;
906: waveform_sig_rx =-1197;
907: waveform_sig_rx =-866;
908: waveform_sig_rx =-939;
909: waveform_sig_rx =-1050;
910: waveform_sig_rx =-1001;
911: waveform_sig_rx =-877;
912: waveform_sig_rx =-940;
913: waveform_sig_rx =-1148;
914: waveform_sig_rx =-785;
915: waveform_sig_rx =-914;
916: waveform_sig_rx =-1113;
917: waveform_sig_rx =-868;
918: waveform_sig_rx =-824;
919: waveform_sig_rx =-1088;
920: waveform_sig_rx =-946;
921: waveform_sig_rx =-737;
922: waveform_sig_rx =-1085;
923: waveform_sig_rx =-985;
924: waveform_sig_rx =-714;
925: waveform_sig_rx =-1009;
926: waveform_sig_rx =-898;
927: waveform_sig_rx =-854;
928: waveform_sig_rx =-975;
929: waveform_sig_rx =-759;
930: waveform_sig_rx =-1027;
931: waveform_sig_rx =-738;
932: waveform_sig_rx =-1065;
933: waveform_sig_rx =-730;
934: waveform_sig_rx =-872;
935: waveform_sig_rx =-1057;
936: waveform_sig_rx =-635;
937: waveform_sig_rx =-946;
938: waveform_sig_rx =-1015;
939: waveform_sig_rx =-574;
940: waveform_sig_rx =-955;
941: waveform_sig_rx =-1003;
942: waveform_sig_rx =-573;
943: waveform_sig_rx =-932;
944: waveform_sig_rx =-929;
945: waveform_sig_rx =-658;
946: waveform_sig_rx =-799;
947: waveform_sig_rx =-960;
948: waveform_sig_rx =-713;
949: waveform_sig_rx =-713;
950: waveform_sig_rx =-852;
951: waveform_sig_rx =-826;
952: waveform_sig_rx =-657;
953: waveform_sig_rx =-752;
954: waveform_sig_rx =-924;
955: waveform_sig_rx =-590;
956: waveform_sig_rx =-741;
957: waveform_sig_rx =-927;
958: waveform_sig_rx =-621;
959: waveform_sig_rx =-622;
960: waveform_sig_rx =-936;
961: waveform_sig_rx =-662;
962: waveform_sig_rx =-588;
963: waveform_sig_rx =-837;
964: waveform_sig_rx =-722;
965: waveform_sig_rx =-593;
966: waveform_sig_rx =-716;
967: waveform_sig_rx =-738;
968: waveform_sig_rx =-667;
969: waveform_sig_rx =-688;
970: waveform_sig_rx =-632;
971: waveform_sig_rx =-734;
972: waveform_sig_rx =-518;
973: waveform_sig_rx =-890;
974: waveform_sig_rx =-417;
975: waveform_sig_rx =-711;
976: waveform_sig_rx =-784;
977: waveform_sig_rx =-370;
978: waveform_sig_rx =-796;
979: waveform_sig_rx =-691;
980: waveform_sig_rx =-376;
981: waveform_sig_rx =-737;
982: waveform_sig_rx =-712;
983: waveform_sig_rx =-367;
984: waveform_sig_rx =-684;
985: waveform_sig_rx =-677;
986: waveform_sig_rx =-427;
987: waveform_sig_rx =-568;
988: waveform_sig_rx =-704;
989: waveform_sig_rx =-479;
990: waveform_sig_rx =-490;
991: waveform_sig_rx =-604;
992: waveform_sig_rx =-622;
993: waveform_sig_rx =-360;
994: waveform_sig_rx =-541;
995: waveform_sig_rx =-701;
996: waveform_sig_rx =-248;
997: waveform_sig_rx =-562;
998: waveform_sig_rx =-648;
999: waveform_sig_rx =-355;
1000: waveform_sig_rx =-472;
1001: waveform_sig_rx =-577;
1002: waveform_sig_rx =-470;
1003: waveform_sig_rx =-354;
1004: waveform_sig_rx =-533;
1005: waveform_sig_rx =-561;
1006: waveform_sig_rx =-260;
1007: waveform_sig_rx =-490;
1008: waveform_sig_rx =-518;
1009: waveform_sig_rx =-344;
1010: waveform_sig_rx =-467;
1011: waveform_sig_rx =-367;
1012: waveform_sig_rx =-410;
1013: waveform_sig_rx =-322;
1014: waveform_sig_rx =-580;
1015: waveform_sig_rx =-139;
1016: waveform_sig_rx =-515;
1017: waveform_sig_rx =-449;
1018: waveform_sig_rx =-119;
1019: waveform_sig_rx =-544;
1020: waveform_sig_rx =-378;
1021: waveform_sig_rx =-145;
1022: waveform_sig_rx =-465;
1023: waveform_sig_rx =-414;
1024: waveform_sig_rx =-126;
1025: waveform_sig_rx =-443;
1026: waveform_sig_rx =-380;
1027: waveform_sig_rx =-198;
1028: waveform_sig_rx =-285;
1029: waveform_sig_rx =-427;
1030: waveform_sig_rx =-237;
1031: waveform_sig_rx =-151;
1032: waveform_sig_rx =-377;
1033: waveform_sig_rx =-349;
1034: waveform_sig_rx =-31;
1035: waveform_sig_rx =-361;
1036: waveform_sig_rx =-330;
1037: waveform_sig_rx =0;
1038: waveform_sig_rx =-322;
1039: waveform_sig_rx =-258;
1040: waveform_sig_rx =-148;
1041: waveform_sig_rx =-124;
1042: waveform_sig_rx =-300;
1043: waveform_sig_rx =-235;
1044: waveform_sig_rx =15;
1045: waveform_sig_rx =-298;
1046: waveform_sig_rx =-243;
1047: waveform_sig_rx =62;
1048: waveform_sig_rx =-283;
1049: waveform_sig_rx =-178;
1050: waveform_sig_rx =-70;
1051: waveform_sig_rx =-211;
1052: waveform_sig_rx =-50;
1053: waveform_sig_rx =-156;
1054: waveform_sig_rx =-46;
1055: waveform_sig_rx =-271;
1056: waveform_sig_rx =126;
1057: waveform_sig_rx =-235;
1058: waveform_sig_rx =-139;
1059: waveform_sig_rx =140;
1060: waveform_sig_rx =-266;
1061: waveform_sig_rx =-52;
1062: waveform_sig_rx =101;
1063: waveform_sig_rx =-166;
1064: waveform_sig_rx =-98;
1065: waveform_sig_rx =117;
1066: waveform_sig_rx =-95;
1067: waveform_sig_rx =-148;
1068: waveform_sig_rx =104;
1069: waveform_sig_rx =52;
1070: waveform_sig_rx =-246;
1071: waveform_sig_rx =137;
1072: waveform_sig_rx =80;
1073: waveform_sig_rx =-148;
1074: waveform_sig_rx =23;
1075: waveform_sig_rx =173;
1076: waveform_sig_rx =-57;
1077: waveform_sig_rx =-11;
1078: waveform_sig_rx =202;
1079: waveform_sig_rx =26;
1080: waveform_sig_rx =-21;
1081: waveform_sig_rx =152;
1082: waveform_sig_rx =199;
1083: waveform_sig_rx =-86;
1084: waveform_sig_rx =97;
1085: waveform_sig_rx =286;
1086: waveform_sig_rx =-59;
1087: waveform_sig_rx =73;
1088: waveform_sig_rx =352;
1089: waveform_sig_rx =-16;
1090: waveform_sig_rx =150;
1091: waveform_sig_rx =210;
1092: waveform_sig_rx =66;
1093: waveform_sig_rx =266;
1094: waveform_sig_rx =124;
1095: waveform_sig_rx =243;
1096: waveform_sig_rx =68;
1097: waveform_sig_rx =382;
1098: waveform_sig_rx =63;
1099: waveform_sig_rx =183;
1100: waveform_sig_rx =377;
1101: waveform_sig_rx =93;
1102: waveform_sig_rx =203;
1103: waveform_sig_rx =403;
1104: waveform_sig_rx =152;
1105: waveform_sig_rx =131;
1106: waveform_sig_rx =481;
1107: waveform_sig_rx =169;
1108: waveform_sig_rx =148;
1109: waveform_sig_rx =455;
1110: waveform_sig_rx =289;
1111: waveform_sig_rx =76;
1112: waveform_sig_rx =464;
1113: waveform_sig_rx =331;
1114: waveform_sig_rx =179;
1115: waveform_sig_rx =343;
1116: waveform_sig_rx =422;
1117: waveform_sig_rx =284;
1118: waveform_sig_rx =261;
1119: waveform_sig_rx =481;
1120: waveform_sig_rx =347;
1121: waveform_sig_rx =225;
1122: waveform_sig_rx =477;
1123: waveform_sig_rx =486;
1124: waveform_sig_rx =159;
1125: waveform_sig_rx =475;
1126: waveform_sig_rx =539;
1127: waveform_sig_rx =216;
1128: waveform_sig_rx =413;
1129: waveform_sig_rx =611;
1130: waveform_sig_rx =276;
1131: waveform_sig_rx =441;
1132: waveform_sig_rx =446;
1133: waveform_sig_rx =375;
1134: waveform_sig_rx =544;
1135: waveform_sig_rx =379;
1136: waveform_sig_rx =535;
1137: waveform_sig_rx =340;
1138: waveform_sig_rx =649;
1139: waveform_sig_rx =369;
1140: waveform_sig_rx =408;
1141: waveform_sig_rx =651;
1142: waveform_sig_rx =377;
1143: waveform_sig_rx =423;
1144: waveform_sig_rx =758;
1145: waveform_sig_rx =381;
1146: waveform_sig_rx =407;
1147: waveform_sig_rx =826;
1148: waveform_sig_rx =360;
1149: waveform_sig_rx =490;
1150: waveform_sig_rx =731;
1151: waveform_sig_rx =509;
1152: waveform_sig_rx =410;
1153: waveform_sig_rx =702;
1154: waveform_sig_rx =590;
1155: waveform_sig_rx =498;
1156: waveform_sig_rx =583;
1157: waveform_sig_rx =720;
1158: waveform_sig_rx =549;
1159: waveform_sig_rx =520;
1160: waveform_sig_rx =789;
1161: waveform_sig_rx =600;
1162: waveform_sig_rx =460;
1163: waveform_sig_rx =805;
1164: waveform_sig_rx =695;
1165: waveform_sig_rx =427;
1166: waveform_sig_rx =772;
1167: waveform_sig_rx =745;
1168: waveform_sig_rx =511;
1169: waveform_sig_rx =692;
1170: waveform_sig_rx =805;
1171: waveform_sig_rx =585;
1172: waveform_sig_rx =689;
1173: waveform_sig_rx =692;
1174: waveform_sig_rx =674;
1175: waveform_sig_rx =746;
1176: waveform_sig_rx =653;
1177: waveform_sig_rx =786;
1178: waveform_sig_rx =559;
1179: waveform_sig_rx =912;
1180: waveform_sig_rx =612;
1181: waveform_sig_rx =663;
1182: waveform_sig_rx =942;
1183: waveform_sig_rx =582;
1184: waveform_sig_rx =691;
1185: waveform_sig_rx =1043;
1186: waveform_sig_rx =526;
1187: waveform_sig_rx =718;
1188: waveform_sig_rx =1045;
1189: waveform_sig_rx =529;
1190: waveform_sig_rx =819;
1191: waveform_sig_rx =885;
1192: waveform_sig_rx =744;
1193: waveform_sig_rx =673;
1194: waveform_sig_rx =882;
1195: waveform_sig_rx =875;
1196: waveform_sig_rx =714;
1197: waveform_sig_rx =777;
1198: waveform_sig_rx =993;
1199: waveform_sig_rx =704;
1200: waveform_sig_rx =750;
1201: waveform_sig_rx =1030;
1202: waveform_sig_rx =763;
1203: waveform_sig_rx =731;
1204: waveform_sig_rx =1009;
1205: waveform_sig_rx =885;
1206: waveform_sig_rx =679;
1207: waveform_sig_rx =985;
1208: waveform_sig_rx =926;
1209: waveform_sig_rx =756;
1210: waveform_sig_rx =875;
1211: waveform_sig_rx =1014;
1212: waveform_sig_rx =794;
1213: waveform_sig_rx =873;
1214: waveform_sig_rx =892;
1215: waveform_sig_rx =894;
1216: waveform_sig_rx =903;
1217: waveform_sig_rx =921;
1218: waveform_sig_rx =969;
1219: waveform_sig_rx =747;
1220: waveform_sig_rx =1199;
1221: waveform_sig_rx =741;
1222: waveform_sig_rx =904;
1223: waveform_sig_rx =1166;
1224: waveform_sig_rx =699;
1225: waveform_sig_rx =988;
1226: waveform_sig_rx =1145;
1227: waveform_sig_rx =708;
1228: waveform_sig_rx =989;
1229: waveform_sig_rx =1131;
1230: waveform_sig_rx =800;
1231: waveform_sig_rx =974;
1232: waveform_sig_rx =1051;
1233: waveform_sig_rx =991;
1234: waveform_sig_rx =814;
1235: waveform_sig_rx =1099;
1236: waveform_sig_rx =1044;
1237: waveform_sig_rx =838;
1238: waveform_sig_rx =1013;
1239: waveform_sig_rx =1175;
1240: waveform_sig_rx =875;
1241: waveform_sig_rx =973;
1242: waveform_sig_rx =1208;
1243: waveform_sig_rx =909;
1244: waveform_sig_rx =930;
1245: waveform_sig_rx =1181;
1246: waveform_sig_rx =1006;
1247: waveform_sig_rx =902;
1248: waveform_sig_rx =1113;
1249: waveform_sig_rx =1111;
1250: waveform_sig_rx =935;
1251: waveform_sig_rx =975;
1252: waveform_sig_rx =1232;
1253: waveform_sig_rx =925;
1254: waveform_sig_rx =1034;
1255: waveform_sig_rx =1111;
1256: waveform_sig_rx =1000;
1257: waveform_sig_rx =1087;
1258: waveform_sig_rx =1103;
1259: waveform_sig_rx =1017;
1260: waveform_sig_rx =967;
1261: waveform_sig_rx =1300;
1262: waveform_sig_rx =815;
1263: waveform_sig_rx =1131;
1264: waveform_sig_rx =1216;
1265: waveform_sig_rx =881;
1266: waveform_sig_rx =1145;
1267: waveform_sig_rx =1237;
1268: waveform_sig_rx =893;
1269: waveform_sig_rx =1106;
1270: waveform_sig_rx =1267;
1271: waveform_sig_rx =933;
1272: waveform_sig_rx =1099;
1273: waveform_sig_rx =1200;
1274: waveform_sig_rx =1099;
1275: waveform_sig_rx =919;
1276: waveform_sig_rx =1264;
1277: waveform_sig_rx =1145;
1278: waveform_sig_rx =954;
1279: waveform_sig_rx =1143;
1280: waveform_sig_rx =1264;
1281: waveform_sig_rx =937;
1282: waveform_sig_rx =1127;
1283: waveform_sig_rx =1244;
1284: waveform_sig_rx =1008;
1285: waveform_sig_rx =1071;
1286: waveform_sig_rx =1219;
1287: waveform_sig_rx =1146;
1288: waveform_sig_rx =973;
1289: waveform_sig_rx =1168;
1290: waveform_sig_rx =1249;
1291: waveform_sig_rx =951;
1292: waveform_sig_rx =1129;
1293: waveform_sig_rx =1353;
1294: waveform_sig_rx =913;
1295: waveform_sig_rx =1205;
1296: waveform_sig_rx =1131;
1297: waveform_sig_rx =1065;
1298: waveform_sig_rx =1207;
1299: waveform_sig_rx =1106;
1300: waveform_sig_rx =1118;
1301: waveform_sig_rx =1089;
1302: waveform_sig_rx =1302;
1303: waveform_sig_rx =954;
1304: waveform_sig_rx =1211;
1305: waveform_sig_rx =1274;
1306: waveform_sig_rx =956;
1307: waveform_sig_rx =1184;
1308: waveform_sig_rx =1293;
1309: waveform_sig_rx =942;
1310: waveform_sig_rx =1169;
1311: waveform_sig_rx =1310;
1312: waveform_sig_rx =1001;
1313: waveform_sig_rx =1119;
1314: waveform_sig_rx =1272;
1315: waveform_sig_rx =1148;
1316: waveform_sig_rx =925;
1317: waveform_sig_rx =1351;
1318: waveform_sig_rx =1147;
1319: waveform_sig_rx =998;
1320: waveform_sig_rx =1249;
1321: waveform_sig_rx =1223;
1322: waveform_sig_rx =1023;
1323: waveform_sig_rx =1155;
1324: waveform_sig_rx =1244;
1325: waveform_sig_rx =1107;
1326: waveform_sig_rx =1013;
1327: waveform_sig_rx =1297;
1328: waveform_sig_rx =1193;
1329: waveform_sig_rx =921;
1330: waveform_sig_rx =1294;
1331: waveform_sig_rx =1214;
1332: waveform_sig_rx =960;
1333: waveform_sig_rx =1234;
1334: waveform_sig_rx =1281;
1335: waveform_sig_rx =964;
1336: waveform_sig_rx =1251;
1337: waveform_sig_rx =1076;
1338: waveform_sig_rx =1149;
1339: waveform_sig_rx =1201;
1340: waveform_sig_rx =1122;
1341: waveform_sig_rx =1155;
1342: waveform_sig_rx =1054;
1343: waveform_sig_rx =1309;
1344: waveform_sig_rx =957;
1345: waveform_sig_rx =1187;
1346: waveform_sig_rx =1255;
1347: waveform_sig_rx =988;
1348: waveform_sig_rx =1182;
1349: waveform_sig_rx =1315;
1350: waveform_sig_rx =963;
1351: waveform_sig_rx =1113;
1352: waveform_sig_rx =1359;
1353: waveform_sig_rx =908;
1354: waveform_sig_rx =1102;
1355: waveform_sig_rx =1316;
1356: waveform_sig_rx =1002;
1357: waveform_sig_rx =1002;
1358: waveform_sig_rx =1322;
1359: waveform_sig_rx =1038;
1360: waveform_sig_rx =1063;
1361: waveform_sig_rx =1128;
1362: waveform_sig_rx =1224;
1363: waveform_sig_rx =1008;
1364: waveform_sig_rx =1057;
1365: waveform_sig_rx =1258;
1366: waveform_sig_rx =1029;
1367: waveform_sig_rx =976;
1368: waveform_sig_rx =1283;
1369: waveform_sig_rx =1090;
1370: waveform_sig_rx =892;
1371: waveform_sig_rx =1265;
1372: waveform_sig_rx =1104;
1373: waveform_sig_rx =895;
1374: waveform_sig_rx =1176;
1375: waveform_sig_rx =1176;
1376: waveform_sig_rx =931;
1377: waveform_sig_rx =1188;
1378: waveform_sig_rx =957;
1379: waveform_sig_rx =1153;
1380: waveform_sig_rx =1059;
1381: waveform_sig_rx =1068;
1382: waveform_sig_rx =1094;
1383: waveform_sig_rx =934;
1384: waveform_sig_rx =1270;
1385: waveform_sig_rx =858;
1386: waveform_sig_rx =1074;
1387: waveform_sig_rx =1229;
1388: waveform_sig_rx =818;
1389: waveform_sig_rx =1110;
1390: waveform_sig_rx =1243;
1391: waveform_sig_rx =775;
1392: waveform_sig_rx =1089;
1393: waveform_sig_rx =1219;
1394: waveform_sig_rx =782;
1395: waveform_sig_rx =1077;
1396: waveform_sig_rx =1169;
1397: waveform_sig_rx =884;
1398: waveform_sig_rx =934;
1399: waveform_sig_rx =1159;
1400: waveform_sig_rx =952;
1401: waveform_sig_rx =963;
1402: waveform_sig_rx =973;
1403: waveform_sig_rx =1175;
1404: waveform_sig_rx =841;
1405: waveform_sig_rx =960;
1406: waveform_sig_rx =1172;
1407: waveform_sig_rx =830;
1408: waveform_sig_rx =898;
1409: waveform_sig_rx =1157;
1410: waveform_sig_rx =907;
1411: waveform_sig_rx =811;
1412: waveform_sig_rx =1122;
1413: waveform_sig_rx =953;
1414: waveform_sig_rx =831;
1415: waveform_sig_rx =1047;
1416: waveform_sig_rx =1020;
1417: waveform_sig_rx =850;
1418: waveform_sig_rx =1009;
1419: waveform_sig_rx =854;
1420: waveform_sig_rx =1034;
1421: waveform_sig_rx =842;
1422: waveform_sig_rx =1004;
1423: waveform_sig_rx =910;
1424: waveform_sig_rx =794;
1425: waveform_sig_rx =1165;
1426: waveform_sig_rx =636;
1427: waveform_sig_rx =997;
1428: waveform_sig_rx =1059;
1429: waveform_sig_rx =615;
1430: waveform_sig_rx =1059;
1431: waveform_sig_rx =997;
1432: waveform_sig_rx =631;
1433: waveform_sig_rx =989;
1434: waveform_sig_rx =1007;
1435: waveform_sig_rx =680;
1436: waveform_sig_rx =937;
1437: waveform_sig_rx =978;
1438: waveform_sig_rx =753;
1439: waveform_sig_rx =788;
1440: waveform_sig_rx =977;
1441: waveform_sig_rx =800;
1442: waveform_sig_rx =768;
1443: waveform_sig_rx =798;
1444: waveform_sig_rx =1029;
1445: waveform_sig_rx =601;
1446: waveform_sig_rx =823;
1447: waveform_sig_rx =1010;
1448: waveform_sig_rx =580;
1449: waveform_sig_rx =811;
1450: waveform_sig_rx =939;
1451: waveform_sig_rx =700;
1452: waveform_sig_rx =718;
1453: waveform_sig_rx =851;
1454: waveform_sig_rx =809;
1455: waveform_sig_rx =632;
1456: waveform_sig_rx =795;
1457: waveform_sig_rx =889;
1458: waveform_sig_rx =573;
1459: waveform_sig_rx =824;
1460: waveform_sig_rx =678;
1461: waveform_sig_rx =760;
1462: waveform_sig_rx =670;
1463: waveform_sig_rx =804;
1464: waveform_sig_rx =634;
1465: waveform_sig_rx =674;
1466: waveform_sig_rx =909;
1467: waveform_sig_rx =402;
1468: waveform_sig_rx =853;
1469: waveform_sig_rx =789;
1470: waveform_sig_rx =428;
1471: waveform_sig_rx =879;
1472: waveform_sig_rx =734;
1473: waveform_sig_rx =431;
1474: waveform_sig_rx =781;
1475: waveform_sig_rx =730;
1476: waveform_sig_rx =497;
1477: waveform_sig_rx =697;
1478: waveform_sig_rx =713;
1479: waveform_sig_rx =565;
1480: waveform_sig_rx =487;
1481: waveform_sig_rx =778;
1482: waveform_sig_rx =605;
1483: waveform_sig_rx =446;
1484: waveform_sig_rx =669;
1485: waveform_sig_rx =736;
1486: waveform_sig_rx =338;
1487: waveform_sig_rx =687;
1488: waveform_sig_rx =671;
1489: waveform_sig_rx =410;
1490: waveform_sig_rx =590;
1491: waveform_sig_rx =635;
1492: waveform_sig_rx =518;
1493: waveform_sig_rx =411;
1494: waveform_sig_rx =624;
1495: waveform_sig_rx =582;
1496: waveform_sig_rx =306;
1497: waveform_sig_rx =594;
1498: waveform_sig_rx =636;
1499: waveform_sig_rx =297;
1500: waveform_sig_rx =606;
1501: waveform_sig_rx =401;
1502: waveform_sig_rx =510;
1503: waveform_sig_rx =450;
1504: waveform_sig_rx =529;
1505: waveform_sig_rx =363;
1506: waveform_sig_rx =474;
1507: waveform_sig_rx =612;
1508: waveform_sig_rx =179;
1509: waveform_sig_rx =629;
1510: waveform_sig_rx =460;
1511: waveform_sig_rx =204;
1512: waveform_sig_rx =611;
1513: waveform_sig_rx =425;
1514: waveform_sig_rx =224;
1515: waveform_sig_rx =467;
1516: waveform_sig_rx =469;
1517: waveform_sig_rx =242;
1518: waveform_sig_rx =367;
1519: waveform_sig_rx =519;
1520: waveform_sig_rx =265;
1521: waveform_sig_rx =191;
1522: waveform_sig_rx =571;
1523: waveform_sig_rx =231;
1524: waveform_sig_rx =210;
1525: waveform_sig_rx =427;
1526: waveform_sig_rx =378;
1527: waveform_sig_rx =127;
1528: waveform_sig_rx =386;
1529: waveform_sig_rx =359;
1530: waveform_sig_rx =168;
1531: waveform_sig_rx =249;
1532: waveform_sig_rx =385;
1533: waveform_sig_rx =244;
1534: waveform_sig_rx =81;
1535: waveform_sig_rx =387;
1536: waveform_sig_rx =281;
1537: waveform_sig_rx =26;
1538: waveform_sig_rx =338;
1539: waveform_sig_rx =316;
1540: waveform_sig_rx =4;
1541: waveform_sig_rx =366;
1542: waveform_sig_rx =81;
1543: waveform_sig_rx =239;
1544: waveform_sig_rx =185;
1545: waveform_sig_rx =209;
1546: waveform_sig_rx =85;
1547: waveform_sig_rx =218;
1548: waveform_sig_rx =243;
1549: waveform_sig_rx =-61;
1550: waveform_sig_rx =308;
1551: waveform_sig_rx =130;
1552: waveform_sig_rx =-19;
1553: waveform_sig_rx =204;
1554: waveform_sig_rx =174;
1555: waveform_sig_rx =-88;
1556: waveform_sig_rx =136;
1557: waveform_sig_rx =213;
1558: waveform_sig_rx =-152;
1559: waveform_sig_rx =85;
1560: waveform_sig_rx =218;
1561: waveform_sig_rx =-129;
1562: waveform_sig_rx =-31;
1563: waveform_sig_rx =239;
1564: waveform_sig_rx =-95;
1565: waveform_sig_rx =-45;
1566: waveform_sig_rx =91;
1567: waveform_sig_rx =82;
1568: waveform_sig_rx =-163;
1569: waveform_sig_rx =34;
1570: waveform_sig_rx =72;
1571: waveform_sig_rx =-141;
1572: waveform_sig_rx =-76;
1573: waveform_sig_rx =117;
1574: waveform_sig_rx =-82;
1575: waveform_sig_rx =-233;
1576: waveform_sig_rx =146;
1577: waveform_sig_rx =-77;
1578: waveform_sig_rx =-260;
1579: waveform_sig_rx =91;
1580: waveform_sig_rx =-53;
1581: waveform_sig_rx =-259;
1582: waveform_sig_rx =43;
1583: waveform_sig_rx =-267;
1584: waveform_sig_rx =-16;
1585: waveform_sig_rx =-195;
1586: waveform_sig_rx =-98;
1587: waveform_sig_rx =-203;
1588: waveform_sig_rx =-147;
1589: waveform_sig_rx =-39;
1590: waveform_sig_rx =-362;
1591: waveform_sig_rx =-56;
1592: waveform_sig_rx =-118;
1593: waveform_sig_rx =-391;
1594: waveform_sig_rx =-81;
1595: waveform_sig_rx =-94;
1596: waveform_sig_rx =-467;
1597: waveform_sig_rx =-114;
1598: waveform_sig_rx =-100;
1599: waveform_sig_rx =-489;
1600: waveform_sig_rx =-150;
1601: waveform_sig_rx =-112;
1602: waveform_sig_rx =-432;
1603: waveform_sig_rx =-271;
1604: waveform_sig_rx =-119;
1605: waveform_sig_rx =-379;
1606: waveform_sig_rx =-321;
1607: waveform_sig_rx =-235;
1608: waveform_sig_rx =-216;
1609: waveform_sig_rx =-460;
1610: waveform_sig_rx =-281;
1611: waveform_sig_rx =-190;
1612: waveform_sig_rx =-476;
1613: waveform_sig_rx =-386;
1614: waveform_sig_rx =-149;
1615: waveform_sig_rx =-480;
1616: waveform_sig_rx =-480;
1617: waveform_sig_rx =-172;
1618: waveform_sig_rx =-457;
1619: waveform_sig_rx =-508;
1620: waveform_sig_rx =-255;
1621: waveform_sig_rx =-396;
1622: waveform_sig_rx =-522;
1623: waveform_sig_rx =-327;
1624: waveform_sig_rx =-533;
1625: waveform_sig_rx =-304;
1626: waveform_sig_rx =-547;
1627: waveform_sig_rx =-353;
1628: waveform_sig_rx =-543;
1629: waveform_sig_rx =-461;
1630: waveform_sig_rx =-323;
1631: waveform_sig_rx =-708;
1632: waveform_sig_rx =-334;
1633: waveform_sig_rx =-397;
1634: waveform_sig_rx =-728;
1635: waveform_sig_rx =-313;
1636: waveform_sig_rx =-400;
1637: waveform_sig_rx =-789;
1638: waveform_sig_rx =-308;
1639: waveform_sig_rx =-471;
1640: waveform_sig_rx =-762;
1641: waveform_sig_rx =-396;
1642: waveform_sig_rx =-492;
1643: waveform_sig_rx =-660;
1644: waveform_sig_rx =-578;
1645: waveform_sig_rx =-428;
1646: waveform_sig_rx =-620;
1647: waveform_sig_rx =-655;
1648: waveform_sig_rx =-501;
1649: waveform_sig_rx =-475;
1650: waveform_sig_rx =-780;
1651: waveform_sig_rx =-516;
1652: waveform_sig_rx =-476;
1653: waveform_sig_rx =-781;
1654: waveform_sig_rx =-622;
1655: waveform_sig_rx =-414;
1656: waveform_sig_rx =-777;
1657: waveform_sig_rx =-714;
1658: waveform_sig_rx =-455;
1659: waveform_sig_rx =-718;
1660: waveform_sig_rx =-745;
1661: waveform_sig_rx =-591;
1662: waveform_sig_rx =-619;
1663: waveform_sig_rx =-804;
1664: waveform_sig_rx =-640;
1665: waveform_sig_rx =-746;
1666: waveform_sig_rx =-628;
1667: waveform_sig_rx =-793;
1668: waveform_sig_rx =-579;
1669: waveform_sig_rx =-864;
1670: waveform_sig_rx =-679;
1671: waveform_sig_rx =-594;
1672: waveform_sig_rx =-1007;
1673: waveform_sig_rx =-546;
1674: waveform_sig_rx =-713;
1675: waveform_sig_rx =-1000;
1676: waveform_sig_rx =-531;
1677: waveform_sig_rx =-750;
1678: waveform_sig_rx =-1017;
1679: waveform_sig_rx =-552;
1680: waveform_sig_rx =-796;
1681: waveform_sig_rx =-941;
1682: waveform_sig_rx =-677;
1683: waveform_sig_rx =-756;
1684: waveform_sig_rx =-887;
1685: waveform_sig_rx =-894;
1686: waveform_sig_rx =-649;
1687: waveform_sig_rx =-883;
1688: waveform_sig_rx =-933;
1689: waveform_sig_rx =-710;
1690: waveform_sig_rx =-762;
1691: waveform_sig_rx =-1036;
1692: waveform_sig_rx =-726;
1693: waveform_sig_rx =-750;
1694: waveform_sig_rx =-1040;
1695: waveform_sig_rx =-821;
1696: waveform_sig_rx =-702;
1697: waveform_sig_rx =-1003;
1698: waveform_sig_rx =-896;
1699: waveform_sig_rx =-761;
1700: waveform_sig_rx =-918;
1701: waveform_sig_rx =-990;
1702: waveform_sig_rx =-849;
1703: waveform_sig_rx =-763;
1704: waveform_sig_rx =-1090;
1705: waveform_sig_rx =-816;
1706: waveform_sig_rx =-931;
1707: waveform_sig_rx =-931;
1708: waveform_sig_rx =-930;
1709: waveform_sig_rx =-830;
1710: waveform_sig_rx =-1118;
1711: waveform_sig_rx =-801;
1712: waveform_sig_rx =-908;
1713: waveform_sig_rx =-1176;
1714: waveform_sig_rx =-739;
1715: waveform_sig_rx =-1014;
1716: waveform_sig_rx =-1124;
1717: waveform_sig_rx =-781;
1718: waveform_sig_rx =-973;
1719: waveform_sig_rx =-1189;
1720: waveform_sig_rx =-770;
1721: waveform_sig_rx =-991;
1722: waveform_sig_rx =-1135;
1723: waveform_sig_rx =-889;
1724: waveform_sig_rx =-935;
1725: waveform_sig_rx =-1082;
1726: waveform_sig_rx =-1101;
1727: waveform_sig_rx =-825;
1728: waveform_sig_rx =-1090;
1729: waveform_sig_rx =-1151;
1730: waveform_sig_rx =-849;
1731: waveform_sig_rx =-1002;
1732: waveform_sig_rx =-1235;
1733: waveform_sig_rx =-871;
1734: waveform_sig_rx =-1027;
1735: waveform_sig_rx =-1156;
1736: waveform_sig_rx =-1028;
1737: waveform_sig_rx =-938;
1738: waveform_sig_rx =-1097;
1739: waveform_sig_rx =-1152;
1740: waveform_sig_rx =-889;
1741: waveform_sig_rx =-1075;
1742: waveform_sig_rx =-1229;
1743: waveform_sig_rx =-904;
1744: waveform_sig_rx =-1030;
1745: waveform_sig_rx =-1254;
1746: waveform_sig_rx =-934;
1747: waveform_sig_rx =-1198;
1748: waveform_sig_rx =-1024;
1749: waveform_sig_rx =-1100;
1750: waveform_sig_rx =-1054;
1751: waveform_sig_rx =-1233;
1752: waveform_sig_rx =-988;
1753: waveform_sig_rx =-1079;
1754: waveform_sig_rx =-1278;
1755: waveform_sig_rx =-915;
1756: waveform_sig_rx =-1146;
1757: waveform_sig_rx =-1270;
1758: waveform_sig_rx =-912;
1759: waveform_sig_rx =-1124;
1760: waveform_sig_rx =-1309;
1761: waveform_sig_rx =-942;
1762: waveform_sig_rx =-1116;
1763: waveform_sig_rx =-1244;
1764: waveform_sig_rx =-1046;
1765: waveform_sig_rx =-1002;
1766: waveform_sig_rx =-1254;
1767: waveform_sig_rx =-1206;
1768: waveform_sig_rx =-893;
1769: waveform_sig_rx =-1290;
1770: waveform_sig_rx =-1210;
1771: waveform_sig_rx =-963;
1772: waveform_sig_rx =-1173;
1773: waveform_sig_rx =-1261;
1774: waveform_sig_rx =-1043;
1775: waveform_sig_rx =-1118;
1776: waveform_sig_rx =-1220;
1777: waveform_sig_rx =-1193;
1778: waveform_sig_rx =-959;
1779: waveform_sig_rx =-1283;
1780: waveform_sig_rx =-1263;
1781: waveform_sig_rx =-923;
1782: waveform_sig_rx =-1248;
1783: waveform_sig_rx =-1253;
1784: waveform_sig_rx =-982;
1785: waveform_sig_rx =-1171;
1786: waveform_sig_rx =-1273;
1787: waveform_sig_rx =-1041;
1788: waveform_sig_rx =-1285;
1789: waveform_sig_rx =-1058;
1790: waveform_sig_rx =-1221;
1791: waveform_sig_rx =-1091;
1792: waveform_sig_rx =-1299;
1793: waveform_sig_rx =-1049;
1794: waveform_sig_rx =-1138;
1795: waveform_sig_rx =-1332;
1796: waveform_sig_rx =-974;
1797: waveform_sig_rx =-1200;
1798: waveform_sig_rx =-1268;
1799: waveform_sig_rx =-991;
1800: waveform_sig_rx =-1150;
1801: waveform_sig_rx =-1354;
1802: waveform_sig_rx =-998;
1803: waveform_sig_rx =-1122;
1804: waveform_sig_rx =-1362;
1805: waveform_sig_rx =-1055;
1806: waveform_sig_rx =-1050;
1807: waveform_sig_rx =-1380;
1808: waveform_sig_rx =-1120;
1809: waveform_sig_rx =-1014;
1810: waveform_sig_rx =-1315;
1811: waveform_sig_rx =-1163;
1812: waveform_sig_rx =-1096;
1813: waveform_sig_rx =-1126;
1814: waveform_sig_rx =-1288;
1815: waveform_sig_rx =-1078;
1816: waveform_sig_rx =-1076;
1817: waveform_sig_rx =-1319;
1818: waveform_sig_rx =-1131;
1819: waveform_sig_rx =-982;
1820: waveform_sig_rx =-1330;
1821: waveform_sig_rx =-1206;
1822: waveform_sig_rx =-965;
1823: waveform_sig_rx =-1260;
1824: waveform_sig_rx =-1267;
1825: waveform_sig_rx =-990;
1826: waveform_sig_rx =-1176;
1827: waveform_sig_rx =-1241;
1828: waveform_sig_rx =-1031;
1829: waveform_sig_rx =-1277;
1830: waveform_sig_rx =-1023;
1831: waveform_sig_rx =-1241;
1832: waveform_sig_rx =-1064;
1833: waveform_sig_rx =-1263;
1834: waveform_sig_rx =-1053;
1835: waveform_sig_rx =-1105;
1836: waveform_sig_rx =-1301;
1837: waveform_sig_rx =-987;
1838: waveform_sig_rx =-1139;
1839: waveform_sig_rx =-1312;
1840: waveform_sig_rx =-931;
1841: waveform_sig_rx =-1137;
1842: waveform_sig_rx =-1369;
1843: waveform_sig_rx =-888;
1844: waveform_sig_rx =-1180;
1845: waveform_sig_rx =-1308;
1846: waveform_sig_rx =-977;
1847: waveform_sig_rx =-1090;
1848: waveform_sig_rx =-1282;
1849: waveform_sig_rx =-1064;
1850: waveform_sig_rx =-1013;
1851: waveform_sig_rx =-1200;
1852: waveform_sig_rx =-1156;
1853: waveform_sig_rx =-1029;
1854: waveform_sig_rx =-1048;
1855: waveform_sig_rx =-1276;
1856: waveform_sig_rx =-973;
1857: waveform_sig_rx =-1033;
1858: waveform_sig_rx =-1271;
1859: waveform_sig_rx =-1036;
1860: waveform_sig_rx =-932;
1861: waveform_sig_rx =-1261;
1862: waveform_sig_rx =-1086;
1863: waveform_sig_rx =-894;
1864: waveform_sig_rx =-1188;
1865: waveform_sig_rx =-1120;
1866: waveform_sig_rx =-925;
1867: waveform_sig_rx =-1095;
1868: waveform_sig_rx =-1112;
1869: waveform_sig_rx =-1015;
1870: waveform_sig_rx =-1137;
1871: waveform_sig_rx =-956;
1872: waveform_sig_rx =-1169;
1873: waveform_sig_rx =-910;
1874: waveform_sig_rx =-1225;
1875: waveform_sig_rx =-933;
1876: waveform_sig_rx =-1009;
1877: waveform_sig_rx =-1255;
1878: waveform_sig_rx =-804;
1879: waveform_sig_rx =-1085;
1880: waveform_sig_rx =-1203;
1881: waveform_sig_rx =-739;
1882: waveform_sig_rx =-1113;
1883: waveform_sig_rx =-1189;
1884: waveform_sig_rx =-774;
1885: waveform_sig_rx =-1096;
1886: waveform_sig_rx =-1129;
1887: waveform_sig_rx =-874;
1888: waveform_sig_rx =-966;
1889: waveform_sig_rx =-1155;
1890: waveform_sig_rx =-950;
1891: waveform_sig_rx =-888;
1892: waveform_sig_rx =-1062;
1893: waveform_sig_rx =-1054;
1894: waveform_sig_rx =-848;
1895: waveform_sig_rx =-945;
1896: waveform_sig_rx =-1172;
1897: waveform_sig_rx =-772;
1898: waveform_sig_rx =-931;
1899: waveform_sig_rx =-1147;
1900: waveform_sig_rx =-830;
1901: waveform_sig_rx =-849;
1902: waveform_sig_rx =-1082;
1903: waveform_sig_rx =-931;
1904: waveform_sig_rx =-817;
1905: waveform_sig_rx =-1003;
1906: waveform_sig_rx =-1017;
1907: waveform_sig_rx =-796;
1908: waveform_sig_rx =-922;
1909: waveform_sig_rx =-1022;
1910: waveform_sig_rx =-851;
1911: waveform_sig_rx =-953;
1912: waveform_sig_rx =-841;
1913: waveform_sig_rx =-963;
1914: waveform_sig_rx =-761;
1915: waveform_sig_rx =-1101;
1916: waveform_sig_rx =-680;
1917: waveform_sig_rx =-916;
1918: waveform_sig_rx =-1053;
1919: waveform_sig_rx =-595;
1920: waveform_sig_rx =-1010;
1921: waveform_sig_rx =-960;
1922: waveform_sig_rx =-595;
1923: waveform_sig_rx =-984;
1924: waveform_sig_rx =-939;
1925: waveform_sig_rx =-623;
1926: waveform_sig_rx =-904;
1927: waveform_sig_rx =-909;
1928: waveform_sig_rx =-713;
1929: waveform_sig_rx =-753;
1930: waveform_sig_rx =-962;
1931: waveform_sig_rx =-785;
1932: waveform_sig_rx =-670;
1933: waveform_sig_rx =-885;
1934: waveform_sig_rx =-879;
1935: waveform_sig_rx =-598;
1936: waveform_sig_rx =-791;
1937: waveform_sig_rx =-933;
1938: waveform_sig_rx =-532;
1939: waveform_sig_rx =-813;
1940: waveform_sig_rx =-858;
1941: waveform_sig_rx =-635;
1942: waveform_sig_rx =-693;
1943: waveform_sig_rx =-821;
1944: waveform_sig_rx =-785;
1945: waveform_sig_rx =-574;
1946: waveform_sig_rx =-782;
1947: waveform_sig_rx =-852;
1948: waveform_sig_rx =-504;
1949: waveform_sig_rx =-764;
1950: waveform_sig_rx =-792;
1951: waveform_sig_rx =-602;
1952: waveform_sig_rx =-783;
1953: waveform_sig_rx =-623;
1954: waveform_sig_rx =-711;
1955: waveform_sig_rx =-586;
1956: waveform_sig_rx =-866;
1957: waveform_sig_rx =-420;
1958: waveform_sig_rx =-749;
1959: waveform_sig_rx =-774;
1960: waveform_sig_rx =-381;
1961: waveform_sig_rx =-833;
1962: waveform_sig_rx =-642;
1963: waveform_sig_rx =-409;
1964: waveform_sig_rx =-738;
1965: waveform_sig_rx =-665;
1966: waveform_sig_rx =-478;
1967: waveform_sig_rx =-627;
1968: waveform_sig_rx =-692;
1969: waveform_sig_rx =-496;
1970: waveform_sig_rx =-485;
1971: waveform_sig_rx =-797;
1972: waveform_sig_rx =-502;
1973: waveform_sig_rx =-439;
1974: waveform_sig_rx =-697;
1975: waveform_sig_rx =-579;
1976: waveform_sig_rx =-376;
1977: waveform_sig_rx =-595;
1978: waveform_sig_rx =-640;
1979: waveform_sig_rx =-331;
1980: waveform_sig_rx =-560;
1981: waveform_sig_rx =-577;
1982: waveform_sig_rx =-450;
1983: waveform_sig_rx =-421;
1984: waveform_sig_rx =-572;
1985: waveform_sig_rx =-536;
1986: waveform_sig_rx =-256;
1987: waveform_sig_rx =-576;
1988: waveform_sig_rx =-571;
1989: waveform_sig_rx =-191;
1990: waveform_sig_rx =-550;
1991: waveform_sig_rx =-489;
1992: waveform_sig_rx =-314;
1993: waveform_sig_rx =-554;
1994: waveform_sig_rx =-296;
1995: waveform_sig_rx =-457;
1996: waveform_sig_rx =-332;
1997: waveform_sig_rx =-543;
1998: waveform_sig_rx =-177;
1999: waveform_sig_rx =-494;
2000: waveform_sig_rx =-443;
2001: waveform_sig_rx =-180;
2002: waveform_sig_rx =-515;
2003: waveform_sig_rx =-375;
2004: waveform_sig_rx =-205;
2005: waveform_sig_rx =-407;
2006: waveform_sig_rx =-456;
2007: waveform_sig_rx =-162;
2008: waveform_sig_rx =-351;
2009: waveform_sig_rx =-473;
2010: waveform_sig_rx =-170;
2011: waveform_sig_rx =-232;
2012: waveform_sig_rx =-536;
2013: waveform_sig_rx =-168;
2014: waveform_sig_rx =-194;
2015: waveform_sig_rx =-433;
2016: waveform_sig_rx =-258;
2017: waveform_sig_rx =-135;
2018: waveform_sig_rx =-304;
2019: waveform_sig_rx =-341;
2020: waveform_sig_rx =-102;
2021: waveform_sig_rx =-249;
2022: waveform_sig_rx =-325;
2023: waveform_sig_rx =-164;
2024: waveform_sig_rx =-64;
2025: waveform_sig_rx =-335;
2026: waveform_sig_rx =-206;
2027: waveform_sig_rx =46;
2028: waveform_sig_rx =-354;
2029: waveform_sig_rx =-233;
2030: waveform_sig_rx =80;
2031: waveform_sig_rx =-310;
2032: waveform_sig_rx =-123;
2033: waveform_sig_rx =-102;
2034: waveform_sig_rx =-255;
2035: waveform_sig_rx =27;
2036: waveform_sig_rx =-234;
2037: waveform_sig_rx =-7;
2038: waveform_sig_rx =-242;
2039: waveform_sig_rx =55;
2040: waveform_sig_rx =-158;
2041: waveform_sig_rx =-181;
2042: waveform_sig_rx =100;
2043: waveform_sig_rx =-205;
2044: waveform_sig_rx =-146;
2045: waveform_sig_rx =145;
2046: waveform_sig_rx =-148;
2047: waveform_sig_rx =-193;
2048: waveform_sig_rx =176;
2049: waveform_sig_rx =-91;
2050: waveform_sig_rx =-177;
2051: waveform_sig_rx =167;
2052: waveform_sig_rx =18;
2053: waveform_sig_rx =-214;
2054: waveform_sig_rx =174;
2055: waveform_sig_rx =46;
2056: waveform_sig_rx =-85;
2057: waveform_sig_rx =35;
2058: waveform_sig_rx =117;
2059: waveform_sig_rx =20;
2060: waveform_sig_rx =-69;
2061: waveform_sig_rx =202;
2062: waveform_sig_rx =86;
2063: waveform_sig_rx =-108;
2064: waveform_sig_rx =185;
2065: waveform_sig_rx =220;
2066: waveform_sig_rx =-132;
2067: waveform_sig_rx =172;
2068: waveform_sig_rx =260;
2069: waveform_sig_rx =-59;
2070: waveform_sig_rx =126;
2071: waveform_sig_rx =284;
2072: waveform_sig_rx =17;
2073: waveform_sig_rx =158;
2074: waveform_sig_rx =153;
2075: waveform_sig_rx =112;
2076: waveform_sig_rx =262;
2077: waveform_sig_rx =73;
2078: waveform_sig_rx =305;
2079: waveform_sig_rx =5;
2080: waveform_sig_rx =378;
2081: waveform_sig_rx =132;
2082: waveform_sig_rx =106;
2083: waveform_sig_rx =417;
2084: waveform_sig_rx =78;
2085: waveform_sig_rx =130;
2086: waveform_sig_rx =497;
2087: waveform_sig_rx =103;
2088: waveform_sig_rx =115;
2089: waveform_sig_rx =561;
2090: waveform_sig_rx =96;
2091: waveform_sig_rx =186;
2092: waveform_sig_rx =457;
2093: waveform_sig_rx =237;
2094: waveform_sig_rx =154;
2095: waveform_sig_rx =414;
2096: waveform_sig_rx =325;
2097: waveform_sig_rx =246;
2098: waveform_sig_rx =253;
2099: waveform_sig_rx =467;
2100: waveform_sig_rx =298;
2101: waveform_sig_rx =188;
2102: waveform_sig_rx =548;
2103: waveform_sig_rx =323;
2104: waveform_sig_rx =192;
2105: waveform_sig_rx =512;
2106: waveform_sig_rx =458;
2107: waveform_sig_rx =190;
2108: waveform_sig_rx =486;
2109: waveform_sig_rx =509;
2110: waveform_sig_rx =246;
2111: waveform_sig_rx =417;
2112: waveform_sig_rx =544;
2113: waveform_sig_rx =354;
2114: waveform_sig_rx =418;
2115: waveform_sig_rx =414;
2116: waveform_sig_rx =451;
2117: waveform_sig_rx =484;
2118: waveform_sig_rx =407;
2119: waveform_sig_rx =572;
2120: waveform_sig_rx =257;
2121: waveform_sig_rx =707;
2122: waveform_sig_rx =366;
2123: waveform_sig_rx =361;
2124: waveform_sig_rx =745;
2125: waveform_sig_rx =298;
2126: waveform_sig_rx =459;
2127: waveform_sig_rx =771;
2128: waveform_sig_rx =304;
2129: waveform_sig_rx =458;
2130: waveform_sig_rx =764;
2131: waveform_sig_rx =367;
2132: waveform_sig_rx =500;
2133: waveform_sig_rx =678;
2134: waveform_sig_rx =543;
2135: waveform_sig_rx =433;
2136: waveform_sig_rx =675;
2137: waveform_sig_rx =645;
2138: waveform_sig_rx =479;
2139: waveform_sig_rx =541;
2140: waveform_sig_rx =778;
2141: waveform_sig_rx =512;
2142: waveform_sig_rx =501;
2143: waveform_sig_rx =834;
2144: waveform_sig_rx =563;
2145: waveform_sig_rx =477;
2146: waveform_sig_rx =794;
2147: waveform_sig_rx =674;
2148: waveform_sig_rx =472;
2149: waveform_sig_rx =732;
2150: waveform_sig_rx =721;
2151: waveform_sig_rx =568;
2152: waveform_sig_rx =633;
2153: waveform_sig_rx =811;
2154: waveform_sig_rx =627;
2155: waveform_sig_rx =612;
2156: waveform_sig_rx =742;
2157: waveform_sig_rx =661;
2158: waveform_sig_rx =693;
2159: waveform_sig_rx =724;
2160: waveform_sig_rx =735;
2161: waveform_sig_rx =569;
2162: waveform_sig_rx =1002;
2163: waveform_sig_rx =522;
2164: waveform_sig_rx =715;
2165: waveform_sig_rx =957;
2166: waveform_sig_rx =534;
2167: waveform_sig_rx =785;
2168: waveform_sig_rx =955;
2169: waveform_sig_rx =598;
2170: waveform_sig_rx =726;
2171: waveform_sig_rx =971;
2172: waveform_sig_rx =626;
2173: waveform_sig_rx =753;
2174: waveform_sig_rx =904;
2175: waveform_sig_rx =805;
2176: waveform_sig_rx =640;
2177: waveform_sig_rx =901;
2178: waveform_sig_rx =890;
2179: waveform_sig_rx =691;
2180: waveform_sig_rx =803;
2181: waveform_sig_rx =1015;
2182: waveform_sig_rx =683;
2183: waveform_sig_rx =781;
2184: waveform_sig_rx =1042;
2185: waveform_sig_rx =745;
2186: waveform_sig_rx =788;
2187: waveform_sig_rx =966;
2188: waveform_sig_rx =896;
2189: waveform_sig_rx =758;
2190: waveform_sig_rx =891;
2191: waveform_sig_rx =1012;
2192: waveform_sig_rx =758;
2193: waveform_sig_rx =819;
2194: waveform_sig_rx =1110;
2195: waveform_sig_rx =757;
2196: waveform_sig_rx =880;
2197: waveform_sig_rx =981;
2198: waveform_sig_rx =826;
2199: waveform_sig_rx =990;
2200: waveform_sig_rx =924;
2201: waveform_sig_rx =928;
2202: waveform_sig_rx =833;
2203: waveform_sig_rx =1135;
2204: waveform_sig_rx =761;
2205: waveform_sig_rx =931;
2206: waveform_sig_rx =1113;
2207: waveform_sig_rx =759;
2208: waveform_sig_rx =968;
2209: waveform_sig_rx =1157;
2210: waveform_sig_rx =786;
2211: waveform_sig_rx =946;
2212: waveform_sig_rx =1157;
2213: waveform_sig_rx =815;
2214: waveform_sig_rx =963;
2215: waveform_sig_rx =1057;
2216: waveform_sig_rx =1024;
2217: waveform_sig_rx =764;
2218: waveform_sig_rx =1106;
2219: waveform_sig_rx =1092;
2220: waveform_sig_rx =790;
2221: waveform_sig_rx =1076;
2222: waveform_sig_rx =1127;
2223: waveform_sig_rx =851;
2224: waveform_sig_rx =1025;
2225: waveform_sig_rx =1100;
2226: waveform_sig_rx =988;
2227: waveform_sig_rx =896;
2228: waveform_sig_rx =1105;
2229: waveform_sig_rx =1125;
2230: waveform_sig_rx =789;
2231: waveform_sig_rx =1126;
2232: waveform_sig_rx =1141;
2233: waveform_sig_rx =850;
2234: waveform_sig_rx =1049;
2235: waveform_sig_rx =1208;
2236: waveform_sig_rx =895;
2237: waveform_sig_rx =1067;
2238: waveform_sig_rx =1086;
2239: waveform_sig_rx =1004;
2240: waveform_sig_rx =1131;
2241: waveform_sig_rx =1035;
2242: waveform_sig_rx =1062;
2243: waveform_sig_rx =978;
2244: waveform_sig_rx =1267;
2245: waveform_sig_rx =896;
2246: waveform_sig_rx =1100;
2247: waveform_sig_rx =1206;
2248: waveform_sig_rx =929;
2249: waveform_sig_rx =1087;
2250: waveform_sig_rx =1233;
2251: waveform_sig_rx =946;
2252: waveform_sig_rx =1038;
2253: waveform_sig_rx =1315;
2254: waveform_sig_rx =965;
2255: waveform_sig_rx =1027;
2256: waveform_sig_rx =1259;
2257: waveform_sig_rx =1074;
2258: waveform_sig_rx =871;
2259: waveform_sig_rx =1309;
2260: waveform_sig_rx =1079;
2261: waveform_sig_rx =974;
2262: waveform_sig_rx =1183;
2263: waveform_sig_rx =1179;
2264: waveform_sig_rx =1050;
2265: waveform_sig_rx =1058;
2266: waveform_sig_rx =1238;
2267: waveform_sig_rx =1122;
2268: waveform_sig_rx =949;
2269: waveform_sig_rx =1283;
2270: waveform_sig_rx =1191;
2271: waveform_sig_rx =904;
2272: waveform_sig_rx =1275;
2273: waveform_sig_rx =1185;
2274: waveform_sig_rx =968;
2275: waveform_sig_rx =1166;
2276: waveform_sig_rx =1285;
2277: waveform_sig_rx =979;
2278: waveform_sig_rx =1157;
2279: waveform_sig_rx =1117;
2280: waveform_sig_rx =1099;
2281: waveform_sig_rx =1208;
2282: waveform_sig_rx =1109;
2283: waveform_sig_rx =1145;
2284: waveform_sig_rx =1059;
2285: waveform_sig_rx =1322;
2286: waveform_sig_rx =993;
2287: waveform_sig_rx =1155;
2288: waveform_sig_rx =1270;
2289: waveform_sig_rx =1009;
2290: waveform_sig_rx =1106;
2291: waveform_sig_rx =1388;
2292: waveform_sig_rx =969;
2293: waveform_sig_rx =1084;
2294: waveform_sig_rx =1415;
2295: waveform_sig_rx =900;
2296: waveform_sig_rx =1144;
2297: waveform_sig_rx =1309;
2298: waveform_sig_rx =1036;
2299: waveform_sig_rx =1026;
2300: waveform_sig_rx =1285;
2301: waveform_sig_rx =1098;
2302: waveform_sig_rx =1062;
2303: waveform_sig_rx =1120;
2304: waveform_sig_rx =1269;
2305: waveform_sig_rx =1031;
2306: waveform_sig_rx =1093;
2307: waveform_sig_rx =1313;
2308: waveform_sig_rx =1082;
2309: waveform_sig_rx =1021;
2310: waveform_sig_rx =1312;
2311: waveform_sig_rx =1167;
2312: waveform_sig_rx =929;
2313: waveform_sig_rx =1311;
2314: waveform_sig_rx =1199;
2315: waveform_sig_rx =982;
2316: waveform_sig_rx =1226;
2317: waveform_sig_rx =1269;
2318: waveform_sig_rx =1019;
2319: waveform_sig_rx =1214;
2320: waveform_sig_rx =1084;
2321: waveform_sig_rx =1184;
2322: waveform_sig_rx =1122;
2323: waveform_sig_rx =1094;
2324: waveform_sig_rx =1189;
2325: waveform_sig_rx =979;
2326: waveform_sig_rx =1362;
2327: waveform_sig_rx =963;
2328: waveform_sig_rx =1120;
2329: waveform_sig_rx =1325;
2330: waveform_sig_rx =890;
2331: waveform_sig_rx =1146;
2332: waveform_sig_rx =1359;
2333: waveform_sig_rx =853;
2334: waveform_sig_rx =1160;
2335: waveform_sig_rx =1334;
2336: waveform_sig_rx =899;
2337: waveform_sig_rx =1171;
2338: waveform_sig_rx =1255;
2339: waveform_sig_rx =1055;
2340: waveform_sig_rx =1010;
2341: waveform_sig_rx =1246;
2342: waveform_sig_rx =1099;
2343: waveform_sig_rx =1031;
2344: waveform_sig_rx =1086;
2345: waveform_sig_rx =1255;
2346: waveform_sig_rx =973;
2347: waveform_sig_rx =1049;
2348: waveform_sig_rx =1302;
2349: waveform_sig_rx =1000;
2350: waveform_sig_rx =1006;
2351: waveform_sig_rx =1300;
2352: waveform_sig_rx =1069;
2353: waveform_sig_rx =959;
2354: waveform_sig_rx =1244;
2355: waveform_sig_rx =1120;
2356: waveform_sig_rx =952;
2357: waveform_sig_rx =1101;
2358: waveform_sig_rx =1202;
2359: waveform_sig_rx =959;
2360: waveform_sig_rx =1087;
2361: waveform_sig_rx =1041;
2362: waveform_sig_rx =1104;
2363: waveform_sig_rx =1028;
2364: waveform_sig_rx =1105;
2365: waveform_sig_rx =1038;
2366: waveform_sig_rx =928;
2367: waveform_sig_rx =1310;
2368: waveform_sig_rx =803;
2369: waveform_sig_rx =1105;
2370: waveform_sig_rx =1227;
2371: waveform_sig_rx =784;
2372: waveform_sig_rx =1180;
2373: waveform_sig_rx =1191;
2374: waveform_sig_rx =792;
2375: waveform_sig_rx =1123;
2376: waveform_sig_rx =1154;
2377: waveform_sig_rx =864;
2378: waveform_sig_rx =1063;
2379: waveform_sig_rx =1138;
2380: waveform_sig_rx =982;
2381: waveform_sig_rx =872;
2382: waveform_sig_rx =1161;
2383: waveform_sig_rx =1003;
2384: waveform_sig_rx =888;
2385: waveform_sig_rx =1020;
2386: waveform_sig_rx =1170;
2387: waveform_sig_rx =813;
2388: waveform_sig_rx =995;
2389: waveform_sig_rx =1179;
2390: waveform_sig_rx =825;
2391: waveform_sig_rx =942;
2392: waveform_sig_rx =1133;
2393: waveform_sig_rx =917;
2394: waveform_sig_rx =864;
2395: waveform_sig_rx =1064;
2396: waveform_sig_rx =1032;
2397: waveform_sig_rx =843;
2398: waveform_sig_rx =935;
2399: waveform_sig_rx =1143;
2400: waveform_sig_rx =785;
2401: waveform_sig_rx =996;
2402: waveform_sig_rx =922;
2403: waveform_sig_rx =935;
2404: waveform_sig_rx =930;
2405: waveform_sig_rx =980;
2406: waveform_sig_rx =867;
2407: waveform_sig_rx =854;
2408: waveform_sig_rx =1137;
2409: waveform_sig_rx =620;
2410: waveform_sig_rx =1037;
2411: waveform_sig_rx =1000;
2412: waveform_sig_rx =644;
2413: waveform_sig_rx =1046;
2414: waveform_sig_rx =958;
2415: waveform_sig_rx =695;
2416: waveform_sig_rx =951;
2417: waveform_sig_rx =987;
2418: waveform_sig_rx =745;
2419: waveform_sig_rx =858;
2420: waveform_sig_rx =981;
2421: waveform_sig_rx =820;
2422: waveform_sig_rx =669;
2423: waveform_sig_rx =1037;
2424: waveform_sig_rx =788;
2425: waveform_sig_rx =714;
2426: waveform_sig_rx =882;
2427: waveform_sig_rx =930;
2428: waveform_sig_rx =628;
2429: waveform_sig_rx =851;
2430: waveform_sig_rx =950;
2431: waveform_sig_rx =665;
2432: waveform_sig_rx =771;
2433: waveform_sig_rx =910;
2434: waveform_sig_rx =776;
2435: waveform_sig_rx =653;
2436: waveform_sig_rx =862;
2437: waveform_sig_rx =865;
2438: waveform_sig_rx =566;
2439: waveform_sig_rx =819;
2440: waveform_sig_rx =941;
2441: waveform_sig_rx =510;
2442: waveform_sig_rx =877;
2443: waveform_sig_rx =667;
2444: waveform_sig_rx =719;
2445: waveform_sig_rx =778;
2446: waveform_sig_rx =734;
2447: waveform_sig_rx =657;
2448: waveform_sig_rx =707;
2449: waveform_sig_rx =853;
2450: waveform_sig_rx =461;
2451: waveform_sig_rx =814;
2452: waveform_sig_rx =737;
2453: waveform_sig_rx =500;
2454: waveform_sig_rx =774;
2455: waveform_sig_rx =761;
2456: waveform_sig_rx =483;
2457: waveform_sig_rx =695;
2458: waveform_sig_rx =804;
2459: waveform_sig_rx =476;
2460: waveform_sig_rx =639;
2461: waveform_sig_rx =792;
2462: waveform_sig_rx =521;
2463: waveform_sig_rx =474;
2464: waveform_sig_rx =828;
2465: waveform_sig_rx =522;
2466: waveform_sig_rx =509;
2467: waveform_sig_rx =653;
2468: waveform_sig_rx =672;
2469: waveform_sig_rx =433;
2470: waveform_sig_rx =629;
2471: waveform_sig_rx =682;
2472: waveform_sig_rx =474;
2473: waveform_sig_rx =512;
2474: waveform_sig_rx =665;
2475: waveform_sig_rx =580;
2476: waveform_sig_rx =343;
2477: waveform_sig_rx =702;
2478: waveform_sig_rx =584;
2479: waveform_sig_rx =282;
2480: waveform_sig_rx =658;
2481: waveform_sig_rx =573;
2482: waveform_sig_rx =320;
2483: waveform_sig_rx =650;
2484: waveform_sig_rx =321;
2485: waveform_sig_rx =547;
2486: waveform_sig_rx =446;
2487: waveform_sig_rx =461;
2488: waveform_sig_rx =445;
2489: waveform_sig_rx =388;
2490: waveform_sig_rx =612;
2491: waveform_sig_rx =221;
2492: waveform_sig_rx =530;
2493: waveform_sig_rx =507;
2494: waveform_sig_rx =213;
2495: waveform_sig_rx =519;
2496: waveform_sig_rx =508;
2497: waveform_sig_rx =199;
2498: waveform_sig_rx =438;
2499: waveform_sig_rx =546;
2500: waveform_sig_rx =167;
2501: waveform_sig_rx =370;
2502: waveform_sig_rx =539;
2503: waveform_sig_rx =197;
2504: waveform_sig_rx =258;
2505: waveform_sig_rx =553;
2506: waveform_sig_rx =213;
2507: waveform_sig_rx =310;
2508: waveform_sig_rx =346;
2509: waveform_sig_rx =406;
2510: waveform_sig_rx =190;
2511: waveform_sig_rx =290;
2512: waveform_sig_rx =441;
2513: waveform_sig_rx =168;
2514: waveform_sig_rx =178;
2515: waveform_sig_rx =488;
2516: waveform_sig_rx =205;
2517: waveform_sig_rx =96;
2518: waveform_sig_rx =453;
2519: waveform_sig_rx =214;
2520: waveform_sig_rx =91;
2521: waveform_sig_rx =347;
2522: waveform_sig_rx =264;
2523: waveform_sig_rx =98;
2524: waveform_sig_rx =293;
2525: waveform_sig_rx =85;
2526: waveform_sig_rx =306;
2527: waveform_sig_rx =122;
2528: waveform_sig_rx =247;
2529: waveform_sig_rx =111;
2530: waveform_sig_rx =94;
2531: waveform_sig_rx =334;
2532: waveform_sig_rx =-110;
2533: waveform_sig_rx =245;
2534: waveform_sig_rx =220;
2535: waveform_sig_rx =-107;
2536: waveform_sig_rx =247;
2537: waveform_sig_rx =223;
2538: waveform_sig_rx =-139;
2539: waveform_sig_rx =176;
2540: waveform_sig_rx =239;
2541: waveform_sig_rx =-172;
2542: waveform_sig_rx =144;
2543: waveform_sig_rx =205;
2544: waveform_sig_rx =-128;
2545: waveform_sig_rx =37;
2546: waveform_sig_rx =153;
2547: waveform_sig_rx =-44;
2548: waveform_sig_rx =-9;
2549: waveform_sig_rx =-18;
2550: waveform_sig_rx =174;
2551: waveform_sig_rx =-211;
2552: waveform_sig_rx =7;
2553: waveform_sig_rx =181;
2554: waveform_sig_rx =-211;
2555: waveform_sig_rx =-18;
2556: waveform_sig_rx =139;
2557: waveform_sig_rx =-148;
2558: waveform_sig_rx =-139;
2559: waveform_sig_rx =83;
2560: waveform_sig_rx =-92;
2561: waveform_sig_rx =-217;
2562: waveform_sig_rx =13;
2563: waveform_sig_rx =-4;
2564: waveform_sig_rx =-235;
2565: waveform_sig_rx =-18;
2566: waveform_sig_rx =-216;
2567: waveform_sig_rx =-23;
2568: waveform_sig_rx =-195;
2569: waveform_sig_rx =-29;
2570: waveform_sig_rx =-217;
2571: waveform_sig_rx =-189;
2572: waveform_sig_rx =56;
2573: waveform_sig_rx =-438;
2574: waveform_sig_rx =-38;
2575: waveform_sig_rx =-68;
2576: waveform_sig_rx =-455;
2577: waveform_sig_rx =22;
2578: waveform_sig_rx =-118;
2579: waveform_sig_rx =-486;
2580: waveform_sig_rx =-27;
2581: waveform_sig_rx =-173;
2582: waveform_sig_rx =-422;
2583: waveform_sig_rx =-151;
2584: waveform_sig_rx =-178;
2585: waveform_sig_rx =-329;
2586: waveform_sig_rx =-347;
2587: waveform_sig_rx =-139;
2588: waveform_sig_rx =-319;
2589: waveform_sig_rx =-403;
2590: waveform_sig_rx =-235;
2591: waveform_sig_rx =-159;
2592: waveform_sig_rx =-530;
2593: waveform_sig_rx =-223;
2594: waveform_sig_rx =-182;
2595: waveform_sig_rx =-538;
2596: waveform_sig_rx =-323;
2597: waveform_sig_rx =-199;
2598: waveform_sig_rx =-468;
2599: waveform_sig_rx =-441;
2600: waveform_sig_rx =-239;
2601: waveform_sig_rx =-390;
2602: waveform_sig_rx =-498;
2603: waveform_sig_rx =-330;
2604: waveform_sig_rx =-263;
2605: waveform_sig_rx =-552;
2606: waveform_sig_rx =-352;
2607: waveform_sig_rx =-461;
2608: waveform_sig_rx =-375;
2609: waveform_sig_rx =-485;
2610: waveform_sig_rx =-326;
2611: waveform_sig_rx =-594;
2612: waveform_sig_rx =-397;
2613: waveform_sig_rx =-317;
2614: waveform_sig_rx =-748;
2615: waveform_sig_rx =-263;
2616: waveform_sig_rx =-463;
2617: waveform_sig_rx =-715;
2618: waveform_sig_rx =-286;
2619: waveform_sig_rx =-485;
2620: waveform_sig_rx =-711;
2621: waveform_sig_rx =-381;
2622: waveform_sig_rx =-481;
2623: waveform_sig_rx =-692;
2624: waveform_sig_rx =-476;
2625: waveform_sig_rx =-465;
2626: waveform_sig_rx =-653;
2627: waveform_sig_rx =-675;
2628: waveform_sig_rx =-386;
2629: waveform_sig_rx =-619;
2630: waveform_sig_rx =-723;
2631: waveform_sig_rx =-472;
2632: waveform_sig_rx =-494;
2633: waveform_sig_rx =-814;
2634: waveform_sig_rx =-454;
2635: waveform_sig_rx =-519;
2636: waveform_sig_rx =-768;
2637: waveform_sig_rx =-587;
2638: waveform_sig_rx =-508;
2639: waveform_sig_rx =-675;
2640: waveform_sig_rx =-723;
2641: waveform_sig_rx =-534;
2642: waveform_sig_rx =-629;
2643: waveform_sig_rx =-821;
2644: waveform_sig_rx =-572;
2645: waveform_sig_rx =-553;
2646: waveform_sig_rx =-885;
2647: waveform_sig_rx =-570;
2648: waveform_sig_rx =-756;
2649: waveform_sig_rx =-697;
2650: waveform_sig_rx =-724;
2651: waveform_sig_rx =-657;
2652: waveform_sig_rx =-856;
2653: waveform_sig_rx =-623;
2654: waveform_sig_rx =-662;
2655: waveform_sig_rx =-941;
2656: waveform_sig_rx =-547;
2657: waveform_sig_rx =-779;
2658: waveform_sig_rx =-897;
2659: waveform_sig_rx =-592;
2660: waveform_sig_rx =-731;
2661: waveform_sig_rx =-965;
2662: waveform_sig_rx =-639;
2663: waveform_sig_rx =-707;
2664: waveform_sig_rx =-953;
2665: waveform_sig_rx =-720;
2666: waveform_sig_rx =-683;
2667: waveform_sig_rx =-900;
2668: waveform_sig_rx =-910;
2669: waveform_sig_rx =-603;
2670: waveform_sig_rx =-912;
2671: waveform_sig_rx =-945;
2672: waveform_sig_rx =-665;
2673: waveform_sig_rx =-829;
2674: waveform_sig_rx =-1002;
2675: waveform_sig_rx =-704;
2676: waveform_sig_rx =-836;
2677: waveform_sig_rx =-926;
2678: waveform_sig_rx =-906;
2679: waveform_sig_rx =-716;
2680: waveform_sig_rx =-901;
2681: waveform_sig_rx =-1050;
2682: waveform_sig_rx =-663;
2683: waveform_sig_rx =-927;
2684: waveform_sig_rx =-1061;
2685: waveform_sig_rx =-723;
2686: waveform_sig_rx =-856;
2687: waveform_sig_rx =-1045;
2688: waveform_sig_rx =-768;
2689: waveform_sig_rx =-1024;
2690: waveform_sig_rx =-848;
2691: waveform_sig_rx =-953;
2692: waveform_sig_rx =-867;
2693: waveform_sig_rx =-1054;
2694: waveform_sig_rx =-852;
2695: waveform_sig_rx =-897;
2696: waveform_sig_rx =-1110;
2697: waveform_sig_rx =-782;
2698: waveform_sig_rx =-991;
2699: waveform_sig_rx =-1091;
2700: waveform_sig_rx =-843;
2701: waveform_sig_rx =-914;
2702: waveform_sig_rx =-1162;
2703: waveform_sig_rx =-872;
2704: waveform_sig_rx =-869;
2705: waveform_sig_rx =-1199;
2706: waveform_sig_rx =-918;
2707: waveform_sig_rx =-853;
2708: waveform_sig_rx =-1197;
2709: waveform_sig_rx =-1029;
2710: waveform_sig_rx =-808;
2711: waveform_sig_rx =-1165;
2712: waveform_sig_rx =-1061;
2713: waveform_sig_rx =-924;
2714: waveform_sig_rx =-1019;
2715: waveform_sig_rx =-1153;
2716: waveform_sig_rx =-968;
2717: waveform_sig_rx =-948;
2718: waveform_sig_rx =-1154;
2719: waveform_sig_rx =-1084;
2720: waveform_sig_rx =-836;
2721: waveform_sig_rx =-1172;
2722: waveform_sig_rx =-1163;
2723: waveform_sig_rx =-843;
2724: waveform_sig_rx =-1137;
2725: waveform_sig_rx =-1192;
2726: waveform_sig_rx =-919;
2727: waveform_sig_rx =-1043;
2728: waveform_sig_rx =-1208;
2729: waveform_sig_rx =-958;
2730: waveform_sig_rx =-1217;
2731: waveform_sig_rx =-997;
2732: waveform_sig_rx =-1139;
2733: waveform_sig_rx =-1045;
2734: waveform_sig_rx =-1176;
2735: waveform_sig_rx =-1028;
2736: waveform_sig_rx =-1041;
2737: waveform_sig_rx =-1250;
2738: waveform_sig_rx =-963;
2739: waveform_sig_rx =-1079;
2740: waveform_sig_rx =-1271;
2741: waveform_sig_rx =-950;
2742: waveform_sig_rx =-1018;
2743: waveform_sig_rx =-1409;
2744: waveform_sig_rx =-908;
2745: waveform_sig_rx =-1059;
2746: waveform_sig_rx =-1365;
2747: waveform_sig_rx =-962;
2748: waveform_sig_rx =-1070;
2749: waveform_sig_rx =-1286;
2750: waveform_sig_rx =-1101;
2751: waveform_sig_rx =-996;
2752: waveform_sig_rx =-1220;
2753: waveform_sig_rx =-1192;
2754: waveform_sig_rx =-1054;
2755: waveform_sig_rx =-1077;
2756: waveform_sig_rx =-1304;
2757: waveform_sig_rx =-1066;
2758: waveform_sig_rx =-1036;
2759: waveform_sig_rx =-1297;
2760: waveform_sig_rx =-1161;
2761: waveform_sig_rx =-948;
2762: waveform_sig_rx =-1305;
2763: waveform_sig_rx =-1206;
2764: waveform_sig_rx =-941;
2765: waveform_sig_rx =-1272;
2766: waveform_sig_rx =-1229;
2767: waveform_sig_rx =-1006;
2768: waveform_sig_rx =-1145;
2769: waveform_sig_rx =-1230;
2770: waveform_sig_rx =-1067;
2771: waveform_sig_rx =-1254;
2772: waveform_sig_rx =-1026;
2773: waveform_sig_rx =-1264;
2774: waveform_sig_rx =-1062;
2775: waveform_sig_rx =-1281;
2776: waveform_sig_rx =-1110;
2777: waveform_sig_rx =-1081;
2778: waveform_sig_rx =-1392;
2779: waveform_sig_rx =-999;
2780: waveform_sig_rx =-1136;
2781: waveform_sig_rx =-1406;
2782: waveform_sig_rx =-931;
2783: waveform_sig_rx =-1160;
2784: waveform_sig_rx =-1422;
2785: waveform_sig_rx =-900;
2786: waveform_sig_rx =-1196;
2787: waveform_sig_rx =-1342;
2788: waveform_sig_rx =-1006;
2789: waveform_sig_rx =-1140;
2790: waveform_sig_rx =-1303;
2791: waveform_sig_rx =-1179;
2792: waveform_sig_rx =-1043;
2793: waveform_sig_rx =-1249;
2794: waveform_sig_rx =-1238;
2795: waveform_sig_rx =-1066;
2796: waveform_sig_rx =-1108;
2797: waveform_sig_rx =-1329;
2798: waveform_sig_rx =-1074;
2799: waveform_sig_rx =-1072;
2800: waveform_sig_rx =-1348;
2801: waveform_sig_rx =-1120;
2802: waveform_sig_rx =-975;
2803: waveform_sig_rx =-1364;
2804: waveform_sig_rx =-1144;
2805: waveform_sig_rx =-1022;
2806: waveform_sig_rx =-1263;
2807: waveform_sig_rx =-1190;
2808: waveform_sig_rx =-1087;
2809: waveform_sig_rx =-1093;
2810: waveform_sig_rx =-1279;
2811: waveform_sig_rx =-1100;
2812: waveform_sig_rx =-1190;
2813: waveform_sig_rx =-1109;
2814: waveform_sig_rx =-1219;
2815: waveform_sig_rx =-1011;
2816: waveform_sig_rx =-1344;
2817: waveform_sig_rx =-1005;
2818: waveform_sig_rx =-1092;
2819: waveform_sig_rx =-1374;
2820: waveform_sig_rx =-902;
2821: waveform_sig_rx =-1188;
2822: waveform_sig_rx =-1324;
2823: waveform_sig_rx =-890;
2824: waveform_sig_rx =-1194;
2825: waveform_sig_rx =-1334;
2826: waveform_sig_rx =-892;
2827: waveform_sig_rx =-1196;
2828: waveform_sig_rx =-1257;
2829: waveform_sig_rx =-1004;
2830: waveform_sig_rx =-1098;
2831: waveform_sig_rx =-1213;
2832: waveform_sig_rx =-1138;
2833: waveform_sig_rx =-971;
2834: waveform_sig_rx =-1191;
2835: waveform_sig_rx =-1220;
2836: waveform_sig_rx =-964;
2837: waveform_sig_rx =-1076;
2838: waveform_sig_rx =-1313;
2839: waveform_sig_rx =-914;
2840: waveform_sig_rx =-1058;
2841: waveform_sig_rx =-1254;
2842: waveform_sig_rx =-996;
2843: waveform_sig_rx =-984;
2844: waveform_sig_rx =-1208;
2845: waveform_sig_rx =-1094;
2846: waveform_sig_rx =-949;
2847: waveform_sig_rx =-1116;
2848: waveform_sig_rx =-1199;
2849: waveform_sig_rx =-955;
2850: waveform_sig_rx =-1016;
2851: waveform_sig_rx =-1223;
2852: waveform_sig_rx =-951;
2853: waveform_sig_rx =-1128;
2854: waveform_sig_rx =-1018;
2855: waveform_sig_rx =-1071;
2856: waveform_sig_rx =-949;
2857: waveform_sig_rx =-1248;
2858: waveform_sig_rx =-843;
2859: waveform_sig_rx =-1070;
2860: waveform_sig_rx =-1225;
2861: waveform_sig_rx =-772;
2862: waveform_sig_rx =-1156;
2863: waveform_sig_rx =-1149;
2864: waveform_sig_rx =-808;
2865: waveform_sig_rx =-1112;
2866: waveform_sig_rx =-1167;
2867: waveform_sig_rx =-837;
2868: waveform_sig_rx =-1052;
2869: waveform_sig_rx =-1125;
2870: waveform_sig_rx =-928;
2871: waveform_sig_rx =-914;
2872: waveform_sig_rx =-1131;
2873: waveform_sig_rx =-1009;
2874: waveform_sig_rx =-819;
2875: waveform_sig_rx =-1086;
2876: waveform_sig_rx =-1070;
2877: waveform_sig_rx =-803;
2878: waveform_sig_rx =-989;
2879: waveform_sig_rx =-1155;
2880: waveform_sig_rx =-766;
2881: waveform_sig_rx =-1014;
2882: waveform_sig_rx =-1086;
2883: waveform_sig_rx =-890;
2884: waveform_sig_rx =-892;
2885: waveform_sig_rx =-1021;
2886: waveform_sig_rx =-1011;
2887: waveform_sig_rx =-790;
2888: waveform_sig_rx =-958;
2889: waveform_sig_rx =-1100;
2890: waveform_sig_rx =-733;
2891: waveform_sig_rx =-924;
2892: waveform_sig_rx =-1062;
2893: waveform_sig_rx =-741;
2894: waveform_sig_rx =-1046;
2895: waveform_sig_rx =-818;
2896: waveform_sig_rx =-918;
2897: waveform_sig_rx =-833;
2898: waveform_sig_rx =-1031;
2899: waveform_sig_rx =-712;
2900: waveform_sig_rx =-936;
2901: waveform_sig_rx =-990;
2902: waveform_sig_rx =-660;
2903: waveform_sig_rx =-986;
2904: waveform_sig_rx =-936;
2905: waveform_sig_rx =-666;
2906: waveform_sig_rx =-902;
2907: waveform_sig_rx =-960;
2908: waveform_sig_rx =-664;
2909: waveform_sig_rx =-829;
2910: waveform_sig_rx =-956;
2911: waveform_sig_rx =-740;
2912: waveform_sig_rx =-714;
2913: waveform_sig_rx =-1022;
2914: waveform_sig_rx =-761;
2915: waveform_sig_rx =-636;
2916: waveform_sig_rx =-973;
2917: waveform_sig_rx =-799;
2918: waveform_sig_rx =-654;
2919: waveform_sig_rx =-841;
2920: waveform_sig_rx =-880;
2921: waveform_sig_rx =-612;
2922: waveform_sig_rx =-761;
2923: waveform_sig_rx =-850;
2924: waveform_sig_rx =-723;
2925: waveform_sig_rx =-629;
2926: waveform_sig_rx =-851;
2927: waveform_sig_rx =-835;
2928: waveform_sig_rx =-498;
2929: waveform_sig_rx =-844;
2930: waveform_sig_rx =-860;
2931: waveform_sig_rx =-460;
2932: waveform_sig_rx =-811;
2933: waveform_sig_rx =-753;
2934: waveform_sig_rx =-561;
2935: waveform_sig_rx =-859;
2936: waveform_sig_rx =-512;
2937: waveform_sig_rx =-746;
2938: waveform_sig_rx =-603;
2939: waveform_sig_rx =-795;
2940: waveform_sig_rx =-537;
2941: waveform_sig_rx =-689;
2942: waveform_sig_rx =-776;
2943: waveform_sig_rx =-459;
2944: waveform_sig_rx =-715;
2945: waveform_sig_rx =-721;
2946: waveform_sig_rx =-401;
2947: waveform_sig_rx =-675;
2948: waveform_sig_rx =-741;
2949: waveform_sig_rx =-426;
2950: waveform_sig_rx =-600;
2951: waveform_sig_rx =-744;
2952: waveform_sig_rx =-460;
2953: waveform_sig_rx =-452;
2954: waveform_sig_rx =-814;
2955: waveform_sig_rx =-437;
2956: waveform_sig_rx =-452;
2957: waveform_sig_rx =-720;
2958: waveform_sig_rx =-487;
2959: waveform_sig_rx =-482;
2960: waveform_sig_rx =-521;
2961: waveform_sig_rx =-651;
2962: waveform_sig_rx =-435;
2963: waveform_sig_rx =-424;
2964: waveform_sig_rx =-684;
2965: waveform_sig_rx =-437;
2966: waveform_sig_rx =-320;
2967: waveform_sig_rx =-692;
2968: waveform_sig_rx =-476;
2969: waveform_sig_rx =-315;
2970: waveform_sig_rx =-612;
2971: waveform_sig_rx =-512;
2972: waveform_sig_rx =-258;
2973: waveform_sig_rx =-527;
2974: waveform_sig_rx =-468;
2975: waveform_sig_rx =-372;
2976: waveform_sig_rx =-537;
2977: waveform_sig_rx =-282;
2978: waveform_sig_rx =-528;
2979: waveform_sig_rx =-291;
2980: waveform_sig_rx =-569;
2981: waveform_sig_rx =-252;
2982: waveform_sig_rx =-401;
2983: waveform_sig_rx =-518;
2984: waveform_sig_rx =-175;
2985: waveform_sig_rx =-444;
2986: waveform_sig_rx =-477;
2987: waveform_sig_rx =-132;
2988: waveform_sig_rx =-404;
2989: waveform_sig_rx =-539;
2990: waveform_sig_rx =-91;
2991: waveform_sig_rx =-379;
2992: waveform_sig_rx =-484;
2993: waveform_sig_rx =-110;
2994: waveform_sig_rx =-293;
2995: waveform_sig_rx =-484;
2996: waveform_sig_rx =-140;
2997: waveform_sig_rx =-263;
2998: waveform_sig_rx =-334;
2999: waveform_sig_rx =-300;
3000: waveform_sig_rx =-194;
3001: waveform_sig_rx =-199;
3002: waveform_sig_rx =-454;
3003: waveform_sig_rx =-39;
3004: waveform_sig_rx =-206;
3005: waveform_sig_rx =-436;
3006: waveform_sig_rx =-76;
3007: waveform_sig_rx =-112;
3008: waveform_sig_rx =-371;
3009: waveform_sig_rx =-167;
3010: waveform_sig_rx =-43;
3011: waveform_sig_rx =-303;
3012: waveform_sig_rx =-239;
3013: waveform_sig_rx =-1;
3014: waveform_sig_rx =-249;
3015: waveform_sig_rx =-180;
3016: waveform_sig_rx =-118;
3017: waveform_sig_rx =-204;
3018: waveform_sig_rx =-27;
3019: waveform_sig_rx =-247;
3020: waveform_sig_rx =18;
3021: waveform_sig_rx =-303;
3022: waveform_sig_rx =57;
3023: waveform_sig_rx =-127;
3024: waveform_sig_rx =-267;
3025: waveform_sig_rx =164;
3026: waveform_sig_rx =-202;
3027: waveform_sig_rx =-210;
3028: waveform_sig_rx =223;
3029: waveform_sig_rx =-221;
3030: waveform_sig_rx =-190;
3031: waveform_sig_rx =222;
3032: waveform_sig_rx =-166;
3033: waveform_sig_rx =-104;
3034: waveform_sig_rx =127;
3035: waveform_sig_rx =-28;
3036: waveform_sig_rx =-151;
3037: waveform_sig_rx =70;
3038: waveform_sig_rx =97;
3039: waveform_sig_rx =-45;
3040: waveform_sig_rx =-64;
3041: waveform_sig_rx =197;
3042: waveform_sig_rx =6;
3043: waveform_sig_rx =-131;
3044: waveform_sig_rx =293;
3045: waveform_sig_rx =18;
3046: waveform_sig_rx =-73;
3047: waveform_sig_rx =200;
3048: waveform_sig_rx =147;
3049: waveform_sig_rx =-67;
3050: waveform_sig_rx =117;
3051: waveform_sig_rx =219;
3052: waveform_sig_rx =-9;
3053: waveform_sig_rx =41;
3054: waveform_sig_rx =276;
3055: waveform_sig_rx =77;
3056: waveform_sig_rx =70;
3057: waveform_sig_rx =153;
3058: waveform_sig_rx =126;
3059: waveform_sig_rx =188;
3060: waveform_sig_rx =114;
3061: waveform_sig_rx =279;
3062: waveform_sig_rx =-59;
3063: waveform_sig_rx =429;
3064: waveform_sig_rx =82;
3065: waveform_sig_rx =82;
3066: waveform_sig_rx =497;
3067: waveform_sig_rx =5;
3068: waveform_sig_rx =195;
3069: waveform_sig_rx =456;
3070: waveform_sig_rx =77;
3071: waveform_sig_rx =194;
3072: waveform_sig_rx =429;
3073: waveform_sig_rx =181;
3074: waveform_sig_rx =185;
3075: waveform_sig_rx =389;
3076: waveform_sig_rx =326;
3077: waveform_sig_rx =91;
3078: waveform_sig_rx =394;
3079: waveform_sig_rx =404;
3080: waveform_sig_rx =208;
3081: waveform_sig_rx =267;
3082: waveform_sig_rx =496;
3083: waveform_sig_rx =259;
3084: waveform_sig_rx =194;
3085: waveform_sig_rx =566;
3086: waveform_sig_rx =278;
3087: waveform_sig_rx =240;
3088: waveform_sig_rx =488;
3089: waveform_sig_rx =394;
3090: waveform_sig_rx =265;
3091: waveform_sig_rx =370;
3092: waveform_sig_rx =511;
3093: waveform_sig_rx =328;
3094: waveform_sig_rx =282;
3095: waveform_sig_rx =637;
3096: waveform_sig_rx =326;
3097: waveform_sig_rx =353;
3098: waveform_sig_rx =529;
3099: waveform_sig_rx =331;
3100: waveform_sig_rx =507;
3101: waveform_sig_rx =423;
3102: waveform_sig_rx =482;
3103: waveform_sig_rx =304;
3104: waveform_sig_rx =707;
3105: waveform_sig_rx =293;
3106: waveform_sig_rx =449;
3107: waveform_sig_rx =698;
3108: waveform_sig_rx =320;
3109: waveform_sig_rx =493;
3110: waveform_sig_rx =693;
3111: waveform_sig_rx =386;
3112: waveform_sig_rx =428;
3113: waveform_sig_rx =727;
3114: waveform_sig_rx =427;
3115: waveform_sig_rx =452;
3116: waveform_sig_rx =653;
3117: waveform_sig_rx =586;
3118: waveform_sig_rx =347;
3119: waveform_sig_rx =655;
3120: waveform_sig_rx =672;
3121: waveform_sig_rx =414;
3122: waveform_sig_rx =567;
3123: waveform_sig_rx =751;
3124: waveform_sig_rx =455;
3125: waveform_sig_rx =541;
3126: waveform_sig_rx =768;
3127: waveform_sig_rx =558;
3128: waveform_sig_rx =542;
3129: waveform_sig_rx =695;
3130: waveform_sig_rx =741;
3131: waveform_sig_rx =494;
3132: waveform_sig_rx =649;
3133: waveform_sig_rx =840;
3134: waveform_sig_rx =502;
3135: waveform_sig_rx =613;
3136: waveform_sig_rx =890;
3137: waveform_sig_rx =524;
3138: waveform_sig_rx =677;
3139: waveform_sig_rx =758;
3140: waveform_sig_rx =587;
3141: waveform_sig_rx =811;
3142: waveform_sig_rx =658;
3143: waveform_sig_rx =742;
3144: waveform_sig_rx =585;
3145: waveform_sig_rx =901;
3146: waveform_sig_rx =569;
3147: waveform_sig_rx =701;
3148: waveform_sig_rx =885;
3149: waveform_sig_rx =582;
3150: waveform_sig_rx =715;
3151: waveform_sig_rx =934;
3152: waveform_sig_rx =642;
3153: waveform_sig_rx =651;
3154: waveform_sig_rx =997;
3155: waveform_sig_rx =671;
3156: waveform_sig_rx =665;
3157: waveform_sig_rx =930;
3158: waveform_sig_rx =796;
3159: waveform_sig_rx =559;
3160: waveform_sig_rx =952;
3161: waveform_sig_rx =845;
3162: waveform_sig_rx =641;
3163: waveform_sig_rx =821;
3164: waveform_sig_rx =922;
3165: waveform_sig_rx =749;
3166: waveform_sig_rx =771;
3167: waveform_sig_rx =954;
3168: waveform_sig_rx =849;
3169: waveform_sig_rx =696;
3170: waveform_sig_rx =924;
3171: waveform_sig_rx =988;
3172: waveform_sig_rx =628;
3173: waveform_sig_rx =954;
3174: waveform_sig_rx =1006;
3175: waveform_sig_rx =682;
3176: waveform_sig_rx =887;
3177: waveform_sig_rx =1048;
3178: waveform_sig_rx =768;
3179: waveform_sig_rx =914;
3180: waveform_sig_rx =924;
3181: waveform_sig_rx =857;
3182: waveform_sig_rx =990;
3183: waveform_sig_rx =857;
3184: waveform_sig_rx =976;
3185: waveform_sig_rx =806;
3186: waveform_sig_rx =1092;
3187: waveform_sig_rx =815;
3188: waveform_sig_rx =901;
3189: waveform_sig_rx =1090;
3190: waveform_sig_rx =827;
3191: waveform_sig_rx =851;
3192: waveform_sig_rx =1166;
3193: waveform_sig_rx =819;
3194: waveform_sig_rx =827;
3195: waveform_sig_rx =1244;
3196: waveform_sig_rx =791;
3197: waveform_sig_rx =904;
3198: waveform_sig_rx =1160;
3199: waveform_sig_rx =897;
3200: waveform_sig_rx =848;
3201: waveform_sig_rx =1140;
3202: waveform_sig_rx =989;
3203: waveform_sig_rx =906;
3204: waveform_sig_rx =979;
3205: waveform_sig_rx =1132;
3206: waveform_sig_rx =921;
3207: waveform_sig_rx =910;
3208: waveform_sig_rx =1165;
3209: waveform_sig_rx =984;
3210: waveform_sig_rx =875;
3211: waveform_sig_rx =1144;
3212: waveform_sig_rx =1116;
3213: waveform_sig_rx =798;
3214: waveform_sig_rx =1154;
3215: waveform_sig_rx =1145;
3216: waveform_sig_rx =855;
3217: waveform_sig_rx =1100;
3218: waveform_sig_rx =1157;
3219: waveform_sig_rx =951;
3220: waveform_sig_rx =1066;
3221: waveform_sig_rx =1010;
3222: waveform_sig_rx =1044;
3223: waveform_sig_rx =1083;
3224: waveform_sig_rx =1001;
3225: waveform_sig_rx =1145;
3226: waveform_sig_rx =868;
3227: waveform_sig_rx =1277;
3228: waveform_sig_rx =953;
3229: waveform_sig_rx =1004;
3230: waveform_sig_rx =1306;
3231: waveform_sig_rx =899;
3232: waveform_sig_rx =1026;
3233: waveform_sig_rx =1356;
3234: waveform_sig_rx =861;
3235: waveform_sig_rx =1028;
3236: waveform_sig_rx =1366;
3237: waveform_sig_rx =860;
3238: waveform_sig_rx =1097;
3239: waveform_sig_rx =1232;
3240: waveform_sig_rx =1021;
3241: waveform_sig_rx =988;
3242: waveform_sig_rx =1209;
3243: waveform_sig_rx =1129;
3244: waveform_sig_rx =1022;
3245: waveform_sig_rx =1078;
3246: waveform_sig_rx =1285;
3247: waveform_sig_rx =1016;
3248: waveform_sig_rx =1046;
3249: waveform_sig_rx =1315;
3250: waveform_sig_rx =1041;
3251: waveform_sig_rx =980;
3252: waveform_sig_rx =1292;
3253: waveform_sig_rx =1127;
3254: waveform_sig_rx =914;
3255: waveform_sig_rx =1283;
3256: waveform_sig_rx =1153;
3257: waveform_sig_rx =1021;
3258: waveform_sig_rx =1158;
3259: waveform_sig_rx =1249;
3260: waveform_sig_rx =1079;
3261: waveform_sig_rx =1098;
3262: waveform_sig_rx =1144;
3263: waveform_sig_rx =1150;
3264: waveform_sig_rx =1134;
3265: waveform_sig_rx =1163;
3266: waveform_sig_rx =1165;
3267: waveform_sig_rx =996;
3268: waveform_sig_rx =1384;
3269: waveform_sig_rx =942;
3270: waveform_sig_rx =1128;
3271: waveform_sig_rx =1331;
3272: waveform_sig_rx =901;
3273: waveform_sig_rx =1156;
3274: waveform_sig_rx =1348;
3275: waveform_sig_rx =897;
3276: waveform_sig_rx =1151;
3277: waveform_sig_rx =1345;
3278: waveform_sig_rx =920;
3279: waveform_sig_rx =1189;
3280: waveform_sig_rx =1244;
3281: waveform_sig_rx =1098;
3282: waveform_sig_rx =1017;
3283: waveform_sig_rx =1232;
3284: waveform_sig_rx =1198;
3285: waveform_sig_rx =1029;
3286: waveform_sig_rx =1125;
3287: waveform_sig_rx =1329;
3288: waveform_sig_rx =992;
3289: waveform_sig_rx =1094;
3290: waveform_sig_rx =1351;
3291: waveform_sig_rx =1022;
3292: waveform_sig_rx =1064;
3293: waveform_sig_rx =1312;
3294: waveform_sig_rx =1126;
3295: waveform_sig_rx =1028;
3296: waveform_sig_rx =1234;
3297: waveform_sig_rx =1206;
3298: waveform_sig_rx =1043;
3299: waveform_sig_rx =1102;
3300: waveform_sig_rx =1318;
3301: waveform_sig_rx =1003;
3302: waveform_sig_rx =1120;
3303: waveform_sig_rx =1175;
3304: waveform_sig_rx =1091;
3305: waveform_sig_rx =1140;
3306: waveform_sig_rx =1163;
3307: waveform_sig_rx =1099;
3308: waveform_sig_rx =1021;
3309: waveform_sig_rx =1376;
3310: waveform_sig_rx =902;
3311: waveform_sig_rx =1189;
3312: waveform_sig_rx =1295;
3313: waveform_sig_rx =907;
3314: waveform_sig_rx =1217;
3315: waveform_sig_rx =1307;
3316: waveform_sig_rx =922;
3317: waveform_sig_rx =1165;
3318: waveform_sig_rx =1294;
3319: waveform_sig_rx =969;
3320: waveform_sig_rx =1158;
3321: waveform_sig_rx =1204;
3322: waveform_sig_rx =1137;
3323: waveform_sig_rx =935;
3324: waveform_sig_rx =1252;
3325: waveform_sig_rx =1168;
3326: waveform_sig_rx =942;
3327: waveform_sig_rx =1144;
3328: waveform_sig_rx =1260;
3329: waveform_sig_rx =928;
3330: waveform_sig_rx =1133;
3331: waveform_sig_rx =1270;
3332: waveform_sig_rx =1003;
3333: waveform_sig_rx =1051;
3334: waveform_sig_rx =1209;
3335: waveform_sig_rx =1107;
3336: waveform_sig_rx =954;
3337: waveform_sig_rx =1182;
3338: waveform_sig_rx =1196;
3339: waveform_sig_rx =950;
3340: waveform_sig_rx =1072;
3341: waveform_sig_rx =1296;
3342: waveform_sig_rx =893;
3343: waveform_sig_rx =1109;
3344: waveform_sig_rx =1111;
3345: waveform_sig_rx =1002;
3346: waveform_sig_rx =1144;
3347: waveform_sig_rx =1084;
3348: waveform_sig_rx =1020;
3349: waveform_sig_rx =1018;
3350: waveform_sig_rx =1239;
3351: waveform_sig_rx =847;
3352: waveform_sig_rx =1159;
3353: waveform_sig_rx =1163;
3354: waveform_sig_rx =871;
3355: waveform_sig_rx =1101;
3356: waveform_sig_rx =1172;
3357: waveform_sig_rx =865;
3358: waveform_sig_rx =1054;
3359: waveform_sig_rx =1206;
3360: waveform_sig_rx =859;
3361: waveform_sig_rx =1022;
3362: waveform_sig_rx =1144;
3363: waveform_sig_rx =1001;
3364: waveform_sig_rx =832;
3365: waveform_sig_rx =1213;
3366: waveform_sig_rx =1010;
3367: waveform_sig_rx =844;
3368: waveform_sig_rx =1083;
3369: waveform_sig_rx =1112;
3370: waveform_sig_rx =828;
3371: waveform_sig_rx =1022;
3372: waveform_sig_rx =1074;
3373: waveform_sig_rx =906;
3374: waveform_sig_rx =907;
3375: waveform_sig_rx =1087;
3376: waveform_sig_rx =1028;
3377: waveform_sig_rx =793;
3378: waveform_sig_rx =1086;
3379: waveform_sig_rx =1084;
3380: waveform_sig_rx =739;
3381: waveform_sig_rx =1017;
3382: waveform_sig_rx =1113;
3383: waveform_sig_rx =729;
3384: waveform_sig_rx =1059;
3385: waveform_sig_rx =871;
3386: waveform_sig_rx =928;
3387: waveform_sig_rx =984;
3388: waveform_sig_rx =897;
3389: waveform_sig_rx =928;
3390: waveform_sig_rx =854;
3391: waveform_sig_rx =1069;
3392: waveform_sig_rx =720;
3393: waveform_sig_rx =951;
3394: waveform_sig_rx =998;
3395: waveform_sig_rx =716;
3396: waveform_sig_rx =946;
3397: waveform_sig_rx =1027;
3398: waveform_sig_rx =694;
3399: waveform_sig_rx =878;
3400: waveform_sig_rx =1062;
3401: waveform_sig_rx =701;
3402: waveform_sig_rx =833;
3403: waveform_sig_rx =1043;
3404: waveform_sig_rx =780;
3405: waveform_sig_rx =672;
3406: waveform_sig_rx =1079;
3407: waveform_sig_rx =754;
3408: waveform_sig_rx =748;
3409: waveform_sig_rx =890;
3410: waveform_sig_rx =890;
3411: waveform_sig_rx =729;
3412: waveform_sig_rx =793;
3413: waveform_sig_rx =944;
3414: waveform_sig_rx =735;
3415: waveform_sig_rx =687;
3416: waveform_sig_rx =963;
3417: waveform_sig_rx =812;
3418: waveform_sig_rx =578;
3419: waveform_sig_rx =964;
3420: waveform_sig_rx =816;
3421: waveform_sig_rx =572;
3422: waveform_sig_rx =879;
3423: waveform_sig_rx =846;
3424: waveform_sig_rx =608;
3425: waveform_sig_rx =844;
3426: waveform_sig_rx =629;
3427: waveform_sig_rx =789;
3428: waveform_sig_rx =725;
3429: waveform_sig_rx =723;
3430: waveform_sig_rx =720;
3431: waveform_sig_rx =623;
3432: waveform_sig_rx =888;
3433: waveform_sig_rx =501;
3434: waveform_sig_rx =765;
3435: waveform_sig_rx =798;
3436: waveform_sig_rx =481;
3437: waveform_sig_rx =733;
3438: waveform_sig_rx =832;
3439: waveform_sig_rx =467;
3440: waveform_sig_rx =650;
3441: waveform_sig_rx =859;
3442: waveform_sig_rx =408;
3443: waveform_sig_rx =647;
3444: waveform_sig_rx =810;
3445: waveform_sig_rx =459;
3446: waveform_sig_rx =554;
3447: waveform_sig_rx =792;
3448: waveform_sig_rx =505;
3449: waveform_sig_rx =582;
3450: waveform_sig_rx =544;
3451: waveform_sig_rx =753;
3452: waveform_sig_rx =463;
3453: waveform_sig_rx =522;
3454: waveform_sig_rx =801;
3455: waveform_sig_rx =400;
3456: waveform_sig_rx =476;
3457: waveform_sig_rx =746;
3458: waveform_sig_rx =469;
3459: waveform_sig_rx =407;
3460: waveform_sig_rx =672;
3461: waveform_sig_rx =550;
3462: waveform_sig_rx =368;
3463: waveform_sig_rx =580;
3464: waveform_sig_rx =625;
3465: waveform_sig_rx =341;
3466: waveform_sig_rx =611;
3467: waveform_sig_rx =392;
3468: waveform_sig_rx =566;
3469: waveform_sig_rx =445;
3470: waveform_sig_rx =471;
3471: waveform_sig_rx =469;
3472: waveform_sig_rx =333;
3473: waveform_sig_rx =672;
3474: waveform_sig_rx =214;
3475: waveform_sig_rx =482;
3476: waveform_sig_rx =610;
3477: waveform_sig_rx =156;
3478: waveform_sig_rx =524;
3479: waveform_sig_rx =592;
3480: waveform_sig_rx =92;
3481: waveform_sig_rx =528;
3482: waveform_sig_rx =501;
3483: waveform_sig_rx =142;
3484: waveform_sig_rx =468;
3485: waveform_sig_rx =426;
3486: waveform_sig_rx =280;
3487: waveform_sig_rx =264;
3488: waveform_sig_rx =474;
3489: waveform_sig_rx =319;
3490: waveform_sig_rx =249;
3491: waveform_sig_rx =305;
3492: waveform_sig_rx =476;
3493: waveform_sig_rx =99;
3494: waveform_sig_rx =307;
3495: waveform_sig_rx =459;
3496: waveform_sig_rx =93;
3497: waveform_sig_rx =251;
3498: waveform_sig_rx =433;
3499: waveform_sig_rx =174;
3500: waveform_sig_rx =157;
3501: waveform_sig_rx =373;
3502: waveform_sig_rx =251;
3503: waveform_sig_rx =106;
3504: waveform_sig_rx =290;
3505: waveform_sig_rx =316;
3506: waveform_sig_rx =68;
3507: waveform_sig_rx =278;
3508: waveform_sig_rx =125;
3509: waveform_sig_rx =270;
3510: waveform_sig_rx =109;
3511: waveform_sig_rx =256;
3512: waveform_sig_rx =114;
3513: waveform_sig_rx =72;
3514: waveform_sig_rx =392;
3515: waveform_sig_rx =-166;
3516: waveform_sig_rx =257;
3517: waveform_sig_rx =254;
3518: waveform_sig_rx =-205;
3519: waveform_sig_rx =337;
3520: waveform_sig_rx =171;
3521: waveform_sig_rx =-150;
3522: waveform_sig_rx =238;
3523: waveform_sig_rx =127;
3524: waveform_sig_rx =-56;
3525: waveform_sig_rx =89;
3526: waveform_sig_rx =154;
3527: waveform_sig_rx =-9;
3528: waveform_sig_rx =-90;
3529: waveform_sig_rx =223;
3530: waveform_sig_rx =-2;
3531: waveform_sig_rx =-76;
3532: waveform_sig_rx =70;
3533: waveform_sig_rx =152;
3534: waveform_sig_rx =-199;
3535: waveform_sig_rx =48;
3536: waveform_sig_rx =148;
3537: waveform_sig_rx =-219;
3538: waveform_sig_rx =-17;
3539: waveform_sig_rx =105;
3540: waveform_sig_rx =-119;
3541: waveform_sig_rx =-114;
3542: waveform_sig_rx =21;
3543: waveform_sig_rx =-13;
3544: waveform_sig_rx =-214;
3545: waveform_sig_rx =-69;
3546: waveform_sig_rx =97;
3547: waveform_sig_rx =-307;
3548: waveform_sig_rx =-12;
3549: waveform_sig_rx =-142;
3550: waveform_sig_rx =-121;
3551: waveform_sig_rx =-135;
3552: waveform_sig_rx =-63;
3553: waveform_sig_rx =-285;
3554: waveform_sig_rx =-110;
3555: waveform_sig_rx =7;
3556: waveform_sig_rx =-456;
3557: waveform_sig_rx =25;
3558: waveform_sig_rx =-169;
3559: waveform_sig_rx =-384;
3560: waveform_sig_rx =2;
3561: waveform_sig_rx =-157;
3562: waveform_sig_rx =-380;
3563: waveform_sig_rx =-111;
3564: waveform_sig_rx =-134;
3565: waveform_sig_rx =-388;
3566: waveform_sig_rx =-219;
3567: waveform_sig_rx =-127;
3568: waveform_sig_rx =-342;
3569: waveform_sig_rx =-388;
3570: waveform_sig_rx =-76;
3571: waveform_sig_rx =-328;
3572: waveform_sig_rx =-407;
3573: waveform_sig_rx =-235;
3574: waveform_sig_rx =-194;
3575: waveform_sig_rx =-547;
3576: waveform_sig_rx =-197;
3577: waveform_sig_rx =-230;
3578: waveform_sig_rx =-467;
3579: waveform_sig_rx =-315;
3580: waveform_sig_rx =-268;
3581: waveform_sig_rx =-347;
3582: waveform_sig_rx =-521;
3583: waveform_sig_rx =-232;
3584: waveform_sig_rx =-287;
3585: waveform_sig_rx =-597;
3586: waveform_sig_rx =-259;
3587: waveform_sig_rx =-275;
3588: waveform_sig_rx =-625;
3589: waveform_sig_rx =-251;
3590: waveform_sig_rx =-527;
3591: waveform_sig_rx =-375;
3592: waveform_sig_rx =-405;
3593: waveform_sig_rx =-406;
3594: waveform_sig_rx =-533;
3595: waveform_sig_rx =-410;
3596: waveform_sig_rx =-364;
3597: waveform_sig_rx =-675;
3598: waveform_sig_rx =-302;
3599: waveform_sig_rx =-471;
3600: waveform_sig_rx =-651;
3601: waveform_sig_rx =-355;
3602: waveform_sig_rx =-419;
3603: waveform_sig_rx =-686;
3604: waveform_sig_rx =-437;
3605: waveform_sig_rx =-384;
3606: waveform_sig_rx =-693;
3607: waveform_sig_rx =-507;
3608: waveform_sig_rx =-369;
3609: waveform_sig_rx =-669;
3610: waveform_sig_rx =-637;
3611: waveform_sig_rx =-314;
3612: waveform_sig_rx =-677;
3613: waveform_sig_rx =-658;
3614: waveform_sig_rx =-479;
3615: waveform_sig_rx =-531;
3616: waveform_sig_rx =-759;
3617: waveform_sig_rx =-535;
3618: waveform_sig_rx =-544;
3619: waveform_sig_rx =-713;
3620: waveform_sig_rx =-670;
3621: waveform_sig_rx =-472;
3622: waveform_sig_rx =-640;
3623: waveform_sig_rx =-823;
3624: waveform_sig_rx =-445;
3625: waveform_sig_rx =-659;
3626: waveform_sig_rx =-854;
3627: waveform_sig_rx =-493;
3628: waveform_sig_rx =-623;
3629: waveform_sig_rx =-818;
3630: waveform_sig_rx =-523;
3631: waveform_sig_rx =-840;
3632: waveform_sig_rx =-589;
3633: waveform_sig_rx =-745;
3634: waveform_sig_rx =-664;
3635: waveform_sig_rx =-760;
3636: waveform_sig_rx =-702;
3637: waveform_sig_rx =-601;
3638: waveform_sig_rx =-922;
3639: waveform_sig_rx =-627;
3640: waveform_sig_rx =-673;
3641: waveform_sig_rx =-938;
3642: waveform_sig_rx =-628;
3643: waveform_sig_rx =-650;
3644: waveform_sig_rx =-992;
3645: waveform_sig_rx =-650;
3646: waveform_sig_rx =-645;
3647: waveform_sig_rx =-1006;
3648: waveform_sig_rx =-698;
3649: waveform_sig_rx =-653;
3650: waveform_sig_rx =-969;
3651: waveform_sig_rx =-836;
3652: waveform_sig_rx =-618;
3653: waveform_sig_rx =-927;
3654: waveform_sig_rx =-866;
3655: waveform_sig_rx =-782;
3656: waveform_sig_rx =-749;
3657: waveform_sig_rx =-984;
3658: waveform_sig_rx =-794;
3659: waveform_sig_rx =-731;
3660: waveform_sig_rx =-982;
3661: waveform_sig_rx =-923;
3662: waveform_sig_rx =-667;
3663: waveform_sig_rx =-971;
3664: waveform_sig_rx =-996;
3665: waveform_sig_rx =-657;
3666: waveform_sig_rx =-943;
3667: waveform_sig_rx =-992;
3668: waveform_sig_rx =-738;
3669: waveform_sig_rx =-869;
3670: waveform_sig_rx =-1006;
3671: waveform_sig_rx =-795;
3672: waveform_sig_rx =-1017;
3673: waveform_sig_rx =-782;
3674: waveform_sig_rx =-1001;
3675: waveform_sig_rx =-818;
3676: waveform_sig_rx =-1018;
3677: waveform_sig_rx =-933;
3678: waveform_sig_rx =-786;
3679: waveform_sig_rx =-1179;
3680: waveform_sig_rx =-806;
3681: waveform_sig_rx =-884;
3682: waveform_sig_rx =-1188;
3683: waveform_sig_rx =-792;
3684: waveform_sig_rx =-896;
3685: waveform_sig_rx =-1246;
3686: waveform_sig_rx =-801;
3687: waveform_sig_rx =-919;
3688: waveform_sig_rx =-1205;
3689: waveform_sig_rx =-868;
3690: waveform_sig_rx =-926;
3691: waveform_sig_rx =-1143;
3692: waveform_sig_rx =-1030;
3693: waveform_sig_rx =-868;
3694: waveform_sig_rx =-1086;
3695: waveform_sig_rx =-1070;
3696: waveform_sig_rx =-961;
3697: waveform_sig_rx =-908;
3698: waveform_sig_rx =-1228;
3699: waveform_sig_rx =-956;
3700: waveform_sig_rx =-888;
3701: waveform_sig_rx =-1199;
3702: waveform_sig_rx =-1027;
3703: waveform_sig_rx =-841;
3704: waveform_sig_rx =-1178;
3705: waveform_sig_rx =-1084;
3706: waveform_sig_rx =-872;
3707: waveform_sig_rx =-1112;
3708: waveform_sig_rx =-1141;
3709: waveform_sig_rx =-994;
3710: waveform_sig_rx =-972;
3711: waveform_sig_rx =-1196;
3712: waveform_sig_rx =-1012;
3713: waveform_sig_rx =-1124;
3714: waveform_sig_rx =-1040;
3715: waveform_sig_rx =-1140;
3716: waveform_sig_rx =-967;
3717: waveform_sig_rx =-1225;
3718: waveform_sig_rx =-1006;
3719: waveform_sig_rx =-1003;
3720: waveform_sig_rx =-1329;
3721: waveform_sig_rx =-908;
3722: waveform_sig_rx =-1087;
3723: waveform_sig_rx =-1305;
3724: waveform_sig_rx =-894;
3725: waveform_sig_rx =-1044;
3726: waveform_sig_rx =-1362;
3727: waveform_sig_rx =-878;
3728: waveform_sig_rx =-1093;
3729: waveform_sig_rx =-1314;
3730: waveform_sig_rx =-962;
3731: waveform_sig_rx =-1092;
3732: waveform_sig_rx =-1210;
3733: waveform_sig_rx =-1176;
3734: waveform_sig_rx =-1011;
3735: waveform_sig_rx =-1161;
3736: waveform_sig_rx =-1278;
3737: waveform_sig_rx =-1007;
3738: waveform_sig_rx =-1031;
3739: waveform_sig_rx =-1361;
3740: waveform_sig_rx =-977;
3741: waveform_sig_rx =-1077;
3742: waveform_sig_rx =-1295;
3743: waveform_sig_rx =-1088;
3744: waveform_sig_rx =-1017;
3745: waveform_sig_rx =-1221;
3746: waveform_sig_rx =-1209;
3747: waveform_sig_rx =-986;
3748: waveform_sig_rx =-1166;
3749: waveform_sig_rx =-1259;
3750: waveform_sig_rx =-1033;
3751: waveform_sig_rx =-1084;
3752: waveform_sig_rx =-1290;
3753: waveform_sig_rx =-1059;
3754: waveform_sig_rx =-1206;
3755: waveform_sig_rx =-1095;
3756: waveform_sig_rx =-1193;
3757: waveform_sig_rx =-1056;
3758: waveform_sig_rx =-1328;
3759: waveform_sig_rx =-1047;
3760: waveform_sig_rx =-1114;
3761: waveform_sig_rx =-1384;
3762: waveform_sig_rx =-935;
3763: waveform_sig_rx =-1196;
3764: waveform_sig_rx =-1337;
3765: waveform_sig_rx =-939;
3766: waveform_sig_rx =-1173;
3767: waveform_sig_rx =-1349;
3768: waveform_sig_rx =-958;
3769: waveform_sig_rx =-1177;
3770: waveform_sig_rx =-1293;
3771: waveform_sig_rx =-1070;
3772: waveform_sig_rx =-1116;
3773: waveform_sig_rx =-1245;
3774: waveform_sig_rx =-1264;
3775: waveform_sig_rx =-971;
3776: waveform_sig_rx =-1252;
3777: waveform_sig_rx =-1301;
3778: waveform_sig_rx =-988;
3779: waveform_sig_rx =-1179;
3780: waveform_sig_rx =-1334;
3781: waveform_sig_rx =-1002;
3782: waveform_sig_rx =-1149;
3783: waveform_sig_rx =-1260;
3784: waveform_sig_rx =-1178;
3785: waveform_sig_rx =-1025;
3786: waveform_sig_rx =-1257;
3787: waveform_sig_rx =-1262;
3788: waveform_sig_rx =-974;
3789: waveform_sig_rx =-1192;
3790: waveform_sig_rx =-1277;
3791: waveform_sig_rx =-1026;
3792: waveform_sig_rx =-1106;
3793: waveform_sig_rx =-1313;
3794: waveform_sig_rx =-1027;
3795: waveform_sig_rx =-1224;
3796: waveform_sig_rx =-1104;
3797: waveform_sig_rx =-1149;
3798: waveform_sig_rx =-1073;
3799: waveform_sig_rx =-1305;
3800: waveform_sig_rx =-979;
3801: waveform_sig_rx =-1153;
3802: waveform_sig_rx =-1294;
3803: waveform_sig_rx =-914;
3804: waveform_sig_rx =-1218;
3805: waveform_sig_rx =-1228;
3806: waveform_sig_rx =-974;
3807: waveform_sig_rx =-1131;
3808: waveform_sig_rx =-1318;
3809: waveform_sig_rx =-1005;
3810: waveform_sig_rx =-1085;
3811: waveform_sig_rx =-1296;
3812: waveform_sig_rx =-1039;
3813: waveform_sig_rx =-1023;
3814: waveform_sig_rx =-1278;
3815: waveform_sig_rx =-1126;
3816: waveform_sig_rx =-944;
3817: waveform_sig_rx =-1228;
3818: waveform_sig_rx =-1164;
3819: waveform_sig_rx =-971;
3820: waveform_sig_rx =-1128;
3821: waveform_sig_rx =-1237;
3822: waveform_sig_rx =-962;
3823: waveform_sig_rx =-1069;
3824: waveform_sig_rx =-1191;
3825: waveform_sig_rx =-1096;
3826: waveform_sig_rx =-930;
3827: waveform_sig_rx =-1167;
3828: waveform_sig_rx =-1175;
3829: waveform_sig_rx =-870;
3830: waveform_sig_rx =-1146;
3831: waveform_sig_rx =-1227;
3832: waveform_sig_rx =-877;
3833: waveform_sig_rx =-1081;
3834: waveform_sig_rx =-1203;
3835: waveform_sig_rx =-918;
3836: waveform_sig_rx =-1228;
3837: waveform_sig_rx =-940;
3838: waveform_sig_rx =-1089;
3839: waveform_sig_rx =-1017;
3840: waveform_sig_rx =-1153;
3841: waveform_sig_rx =-954;
3842: waveform_sig_rx =-1035;
3843: waveform_sig_rx =-1166;
3844: waveform_sig_rx =-855;
3845: waveform_sig_rx =-1074;
3846: waveform_sig_rx =-1181;
3847: waveform_sig_rx =-845;
3848: waveform_sig_rx =-1004;
3849: waveform_sig_rx =-1226;
3850: waveform_sig_rx =-824;
3851: waveform_sig_rx =-993;
3852: waveform_sig_rx =-1185;
3853: waveform_sig_rx =-878;
3854: waveform_sig_rx =-901;
3855: waveform_sig_rx =-1177;
3856: waveform_sig_rx =-962;
3857: waveform_sig_rx =-824;
3858: waveform_sig_rx =-1129;
3859: waveform_sig_rx =-1010;
3860: waveform_sig_rx =-874;
3861: waveform_sig_rx =-968;
3862: waveform_sig_rx =-1074;
3863: waveform_sig_rx =-892;
3864: waveform_sig_rx =-888;
3865: waveform_sig_rx =-1081;
3866: waveform_sig_rx =-975;
3867: waveform_sig_rx =-753;
3868: waveform_sig_rx =-1103;
3869: waveform_sig_rx =-995;
3870: waveform_sig_rx =-717;
3871: waveform_sig_rx =-1070;
3872: waveform_sig_rx =-999;
3873: waveform_sig_rx =-755;
3874: waveform_sig_rx =-959;
3875: waveform_sig_rx =-978;
3876: waveform_sig_rx =-814;
3877: waveform_sig_rx =-1022;
3878: waveform_sig_rx =-758;
3879: waveform_sig_rx =-997;
3880: waveform_sig_rx =-791;
3881: waveform_sig_rx =-1015;
3882: waveform_sig_rx =-775;
3883: waveform_sig_rx =-819;
3884: waveform_sig_rx =-1040;
3885: waveform_sig_rx =-672;
3886: waveform_sig_rx =-875;
3887: waveform_sig_rx =-1024;
3888: waveform_sig_rx =-630;
3889: waveform_sig_rx =-848;
3890: waveform_sig_rx =-1047;
3891: waveform_sig_rx =-589;
3892: waveform_sig_rx =-846;
3893: waveform_sig_rx =-1009;
3894: waveform_sig_rx =-647;
3895: waveform_sig_rx =-752;
3896: waveform_sig_rx =-982;
3897: waveform_sig_rx =-712;
3898: waveform_sig_rx =-710;
3899: waveform_sig_rx =-883;
3900: waveform_sig_rx =-804;
3901: waveform_sig_rx =-728;
3902: waveform_sig_rx =-718;
3903: waveform_sig_rx =-943;
3904: waveform_sig_rx =-642;
3905: waveform_sig_rx =-656;
3906: waveform_sig_rx =-968;
3907: waveform_sig_rx =-670;
3908: waveform_sig_rx =-597;
3909: waveform_sig_rx =-935;
3910: waveform_sig_rx =-708;
3911: waveform_sig_rx =-555;
3912: waveform_sig_rx =-825;
3913: waveform_sig_rx =-772;
3914: waveform_sig_rx =-570;
3915: waveform_sig_rx =-727;
3916: waveform_sig_rx =-753;
3917: waveform_sig_rx =-616;
3918: waveform_sig_rx =-775;
3919: waveform_sig_rx =-562;
3920: waveform_sig_rx =-771;
3921: waveform_sig_rx =-545;
3922: waveform_sig_rx =-826;
3923: waveform_sig_rx =-544;
3924: waveform_sig_rx =-613;
3925: waveform_sig_rx =-830;
3926: waveform_sig_rx =-434;
3927: waveform_sig_rx =-674;
3928: waveform_sig_rx =-833;
3929: waveform_sig_rx =-359;
3930: waveform_sig_rx =-689;
3931: waveform_sig_rx =-806;
3932: waveform_sig_rx =-324;
3933: waveform_sig_rx =-684;
3934: waveform_sig_rx =-711;
3935: waveform_sig_rx =-418;
3936: waveform_sig_rx =-562;
3937: waveform_sig_rx =-702;
3938: waveform_sig_rx =-518;
3939: waveform_sig_rx =-475;
3940: waveform_sig_rx =-625;
3941: waveform_sig_rx =-626;
3942: waveform_sig_rx =-412;
3943: waveform_sig_rx =-510;
3944: waveform_sig_rx =-712;
3945: waveform_sig_rx =-338;
3946: waveform_sig_rx =-501;
3947: waveform_sig_rx =-677;
3948: waveform_sig_rx =-404;
3949: waveform_sig_rx =-394;
3950: waveform_sig_rx =-636;
3951: waveform_sig_rx =-483;
3952: waveform_sig_rx =-331;
3953: waveform_sig_rx =-563;
3954: waveform_sig_rx =-551;
3955: waveform_sig_rx =-319;
3956: waveform_sig_rx =-461;
3957: waveform_sig_rx =-519;
3958: waveform_sig_rx =-385;
3959: waveform_sig_rx =-475;
3960: waveform_sig_rx =-321;
3961: waveform_sig_rx =-505;
3962: waveform_sig_rx =-252;
3963: waveform_sig_rx =-604;
3964: waveform_sig_rx =-201;
3965: waveform_sig_rx =-402;
3966: waveform_sig_rx =-578;
3967: waveform_sig_rx =-95;
3968: waveform_sig_rx =-514;
3969: waveform_sig_rx =-472;
3970: waveform_sig_rx =-80;
3971: waveform_sig_rx =-483;
3972: waveform_sig_rx =-425;
3973: waveform_sig_rx =-132;
3974: waveform_sig_rx =-397;
3975: waveform_sig_rx =-412;
3976: waveform_sig_rx =-218;
3977: waveform_sig_rx =-241;
3978: waveform_sig_rx =-471;
3979: waveform_sig_rx =-232;
3980: waveform_sig_rx =-158;
3981: waveform_sig_rx =-385;
3982: waveform_sig_rx =-324;
3983: waveform_sig_rx =-135;
3984: waveform_sig_rx =-243;
3985: waveform_sig_rx =-430;
3986: waveform_sig_rx =-39;
3987: waveform_sig_rx =-235;
3988: waveform_sig_rx =-383;
3989: waveform_sig_rx =-93;
3990: waveform_sig_rx =-147;
3991: waveform_sig_rx =-309;
3992: waveform_sig_rx =-185;
3993: waveform_sig_rx =-58;
3994: waveform_sig_rx =-221;
3995: waveform_sig_rx =-293;
3996: waveform_sig_rx =30;
3997: waveform_sig_rx =-196;
3998: waveform_sig_rx =-279;
3999: waveform_sig_rx =-42;
4000: waveform_sig_rx =-230;
4001: waveform_sig_rx =-53;
4002: waveform_sig_rx =-154;
4003: waveform_sig_rx =-37;
4004: waveform_sig_rx =-311;
4005: waveform_sig_rx =113;
4006: waveform_sig_rx =-193;
4007: waveform_sig_rx =-218;
4008: waveform_sig_rx =176;
4009: waveform_sig_rx =-230;
4010: waveform_sig_rx =-98;
4011: waveform_sig_rx =149;
4012: waveform_sig_rx =-165;
4013: waveform_sig_rx =-134;
4014: waveform_sig_rx =147;
4015: waveform_sig_rx =-78;
4016: waveform_sig_rx =-139;
4017: waveform_sig_rx =80;
4018: waveform_sig_rx =72;
4019: waveform_sig_rx =-191;
4020: waveform_sig_rx =74;
4021: waveform_sig_rx =138;
4022: waveform_sig_rx =-110;
4023: waveform_sig_rx =-23;
4024: waveform_sig_rx =164;
4025: waveform_sig_rx =-4;
4026: waveform_sig_rx =-101;
4027: waveform_sig_rx =265;
4028: waveform_sig_rx =17;
4029: waveform_sig_rx =-34;
4030: waveform_sig_rx =167;
4031: waveform_sig_rx =137;
4032: waveform_sig_rx =16;
4033: waveform_sig_rx =29;
4034: waveform_sig_rx =287;
4035: waveform_sig_rx =18;
4036: waveform_sig_rx =-29;
4037: waveform_sig_rx =376;
4038: waveform_sig_rx =14;
4039: waveform_sig_rx =77;
4040: waveform_sig_rx =265;
4041: waveform_sig_rx =20;
4042: waveform_sig_rx =289;
4043: waveform_sig_rx =95;
4044: waveform_sig_rx =245;
4045: waveform_sig_rx =39;
4046: waveform_sig_rx =382;
4047: waveform_sig_rx =132;
4048: waveform_sig_rx =110;
4049: waveform_sig_rx =429;
4050: waveform_sig_rx =86;
4051: waveform_sig_rx =155;
4052: waveform_sig_rx =439;
4053: waveform_sig_rx =120;
4054: waveform_sig_rx =153;
4055: waveform_sig_rx =430;
4056: waveform_sig_rx =211;
4057: waveform_sig_rx =151;
4058: waveform_sig_rx =374;
4059: waveform_sig_rx =391;
4060: waveform_sig_rx =52;
4061: waveform_sig_rx =406;
4062: waveform_sig_rx =398;
4063: waveform_sig_rx =174;
4064: waveform_sig_rx =332;
4065: waveform_sig_rx =429;
4066: waveform_sig_rx =307;
4067: waveform_sig_rx =231;
4068: waveform_sig_rx =498;
4069: waveform_sig_rx =371;
4070: waveform_sig_rx =227;
4071: waveform_sig_rx =439;
4072: waveform_sig_rx =497;
4073: waveform_sig_rx =229;
4074: waveform_sig_rx =377;
4075: waveform_sig_rx =588;
4076: waveform_sig_rx =255;
4077: waveform_sig_rx =340;
4078: waveform_sig_rx =627;
4079: waveform_sig_rx =283;
4080: waveform_sig_rx =421;
4081: waveform_sig_rx =480;
4082: waveform_sig_rx =337;
4083: waveform_sig_rx =564;
4084: waveform_sig_rx =357;
4085: waveform_sig_rx =544;
4086: waveform_sig_rx =286;
4087: waveform_sig_rx =628;
4088: waveform_sig_rx =383;
4089: waveform_sig_rx =368;
4090: waveform_sig_rx =678;
4091: waveform_sig_rx =371;
4092: waveform_sig_rx =426;
4093: waveform_sig_rx =730;
4094: waveform_sig_rx =417;
4095: waveform_sig_rx =393;
4096: waveform_sig_rx =758;
4097: waveform_sig_rx =462;
4098: waveform_sig_rx =400;
4099: waveform_sig_rx =719;
4100: waveform_sig_rx =585;
4101: waveform_sig_rx =353;
4102: waveform_sig_rx =713;
4103: waveform_sig_rx =631;
4104: waveform_sig_rx =486;
4105: waveform_sig_rx =602;
4106: waveform_sig_rx =726;
4107: waveform_sig_rx =587;
4108: waveform_sig_rx =503;
4109: waveform_sig_rx =764;
4110: waveform_sig_rx =643;
4111: waveform_sig_rx =468;
4112: waveform_sig_rx =743;
4113: waveform_sig_rx =767;
4114: waveform_sig_rx =436;
4115: waveform_sig_rx =691;
4116: waveform_sig_rx =807;
4117: waveform_sig_rx =474;
4118: waveform_sig_rx =645;
4119: waveform_sig_rx =822;
4120: waveform_sig_rx =574;
4121: waveform_sig_rx =695;
4122: waveform_sig_rx =692;
4123: waveform_sig_rx =653;
4124: waveform_sig_rx =771;
4125: waveform_sig_rx =596;
4126: waveform_sig_rx =829;
4127: waveform_sig_rx =541;
4128: waveform_sig_rx =916;
4129: waveform_sig_rx =649;
4130: waveform_sig_rx =620;
4131: waveform_sig_rx =955;
4132: waveform_sig_rx =603;
4133: waveform_sig_rx =661;
4134: waveform_sig_rx =977;
4135: waveform_sig_rx =613;
4136: waveform_sig_rx =640;
4137: waveform_sig_rx =1030;
4138: waveform_sig_rx =653;
4139: waveform_sig_rx =689;
4140: waveform_sig_rx =961;
4141: waveform_sig_rx =770;
4142: waveform_sig_rx =626;
4143: waveform_sig_rx =936;
4144: waveform_sig_rx =836;
4145: waveform_sig_rx =738;
4146: waveform_sig_rx =769;
4147: waveform_sig_rx =945;
4148: waveform_sig_rx =784;
4149: waveform_sig_rx =669;
4150: waveform_sig_rx =1022;
4151: waveform_sig_rx =815;
4152: waveform_sig_rx =670;
4153: waveform_sig_rx =1006;
4154: waveform_sig_rx =914;
4155: waveform_sig_rx =654;
4156: waveform_sig_rx =950;
4157: waveform_sig_rx =960;
4158: waveform_sig_rx =758;
4159: waveform_sig_rx =853;
4160: waveform_sig_rx =1011;
4161: waveform_sig_rx =828;
4162: waveform_sig_rx =865;
4163: waveform_sig_rx =907;
4164: waveform_sig_rx =893;
4165: waveform_sig_rx =934;
4166: waveform_sig_rx =880;
4167: waveform_sig_rx =989;
4168: waveform_sig_rx =724;
4169: waveform_sig_rx =1161;
4170: waveform_sig_rx =789;
4171: waveform_sig_rx =843;
4172: waveform_sig_rx =1169;
4173: waveform_sig_rx =766;
4174: waveform_sig_rx =901;
4175: waveform_sig_rx =1199;
4176: waveform_sig_rx =774;
4177: waveform_sig_rx =884;
4178: waveform_sig_rx =1222;
4179: waveform_sig_rx =773;
4180: waveform_sig_rx =937;
4181: waveform_sig_rx =1116;
4182: waveform_sig_rx =936;
4183: waveform_sig_rx =860;
4184: waveform_sig_rx =1054;
4185: waveform_sig_rx =1077;
4186: waveform_sig_rx =918;
4187: waveform_sig_rx =939;
4188: waveform_sig_rx =1216;
4189: waveform_sig_rx =894;
4190: waveform_sig_rx =896;
4191: waveform_sig_rx =1245;
4192: waveform_sig_rx =925;
4193: waveform_sig_rx =927;
4194: waveform_sig_rx =1162;
4195: waveform_sig_rx =1065;
4196: waveform_sig_rx =882;
4197: waveform_sig_rx =1084;
4198: waveform_sig_rx =1148;
4199: waveform_sig_rx =910;
4200: waveform_sig_rx =1020;
4201: waveform_sig_rx =1220;
4202: waveform_sig_rx =946;
4203: waveform_sig_rx =1051;
4204: waveform_sig_rx =1088;
4205: waveform_sig_rx =1023;
4206: waveform_sig_rx =1091;
4207: waveform_sig_rx =1053;
4208: waveform_sig_rx =1112;
4209: waveform_sig_rx =896;
4210: waveform_sig_rx =1314;
4211: waveform_sig_rx =900;
4212: waveform_sig_rx =1017;
4213: waveform_sig_rx =1307;
4214: waveform_sig_rx =859;
4215: waveform_sig_rx =1097;
4216: waveform_sig_rx =1302;
4217: waveform_sig_rx =882;
4218: waveform_sig_rx =1077;
4219: waveform_sig_rx =1275;
4220: waveform_sig_rx =939;
4221: waveform_sig_rx =1084;
4222: waveform_sig_rx =1155;
4223: waveform_sig_rx =1125;
4224: waveform_sig_rx =906;
4225: waveform_sig_rx =1179;
4226: waveform_sig_rx =1207;
4227: waveform_sig_rx =930;
4228: waveform_sig_rx =1121;
4229: waveform_sig_rx =1290;
4230: waveform_sig_rx =940;
4231: waveform_sig_rx =1099;
4232: waveform_sig_rx =1252;
4233: waveform_sig_rx =1057;
4234: waveform_sig_rx =1031;
4235: waveform_sig_rx =1209;
4236: waveform_sig_rx =1191;
4237: waveform_sig_rx =937;
4238: waveform_sig_rx =1185;
4239: waveform_sig_rx =1213;
4240: waveform_sig_rx =1002;
4241: waveform_sig_rx =1105;
4242: waveform_sig_rx =1303;
4243: waveform_sig_rx =1041;
4244: waveform_sig_rx =1107;
4245: waveform_sig_rx =1198;
4246: waveform_sig_rx =1100;
4247: waveform_sig_rx =1147;
4248: waveform_sig_rx =1154;
4249: waveform_sig_rx =1123;
4250: waveform_sig_rx =1023;
4251: waveform_sig_rx =1392;
4252: waveform_sig_rx =928;
4253: waveform_sig_rx =1178;
4254: waveform_sig_rx =1288;
4255: waveform_sig_rx =958;
4256: waveform_sig_rx =1189;
4257: waveform_sig_rx =1283;
4258: waveform_sig_rx =1024;
4259: waveform_sig_rx =1094;
4260: waveform_sig_rx =1344;
4261: waveform_sig_rx =1015;
4262: waveform_sig_rx =1077;
4263: waveform_sig_rx =1284;
4264: waveform_sig_rx =1149;
4265: waveform_sig_rx =956;
4266: waveform_sig_rx =1307;
4267: waveform_sig_rx =1205;
4268: waveform_sig_rx =1007;
4269: waveform_sig_rx =1180;
4270: waveform_sig_rx =1283;
4271: waveform_sig_rx =1014;
4272: waveform_sig_rx =1128;
4273: waveform_sig_rx =1277;
4274: waveform_sig_rx =1080;
4275: waveform_sig_rx =1058;
4276: waveform_sig_rx =1234;
4277: waveform_sig_rx =1211;
4278: waveform_sig_rx =967;
4279: waveform_sig_rx =1218;
4280: waveform_sig_rx =1261;
4281: waveform_sig_rx =975;
4282: waveform_sig_rx =1138;
4283: waveform_sig_rx =1328;
4284: waveform_sig_rx =973;
4285: waveform_sig_rx =1146;
4286: waveform_sig_rx =1156;
4287: waveform_sig_rx =1049;
4288: waveform_sig_rx =1216;
4289: waveform_sig_rx =1124;
4290: waveform_sig_rx =1129;
4291: waveform_sig_rx =1073;
4292: waveform_sig_rx =1332;
4293: waveform_sig_rx =971;
4294: waveform_sig_rx =1166;
4295: waveform_sig_rx =1248;
4296: waveform_sig_rx =1011;
4297: waveform_sig_rx =1118;
4298: waveform_sig_rx =1335;
4299: waveform_sig_rx =989;
4300: waveform_sig_rx =1060;
4301: waveform_sig_rx =1375;
4302: waveform_sig_rx =930;
4303: waveform_sig_rx =1105;
4304: waveform_sig_rx =1256;
4305: waveform_sig_rx =1079;
4306: waveform_sig_rx =964;
4307: waveform_sig_rx =1242;
4308: waveform_sig_rx =1138;
4309: waveform_sig_rx =978;
4310: waveform_sig_rx =1147;
4311: waveform_sig_rx =1233;
4312: waveform_sig_rx =958;
4313: waveform_sig_rx =1106;
4314: waveform_sig_rx =1194;
4315: waveform_sig_rx =1070;
4316: waveform_sig_rx =992;
4317: waveform_sig_rx =1211;
4318: waveform_sig_rx =1192;
4319: waveform_sig_rx =837;
4320: waveform_sig_rx =1238;
4321: waveform_sig_rx =1192;
4322: waveform_sig_rx =876;
4323: waveform_sig_rx =1181;
4324: waveform_sig_rx =1201;
4325: waveform_sig_rx =943;
4326: waveform_sig_rx =1135;
4327: waveform_sig_rx =1018;
4328: waveform_sig_rx =1074;
4329: waveform_sig_rx =1098;
4330: waveform_sig_rx =1032;
4331: waveform_sig_rx =1087;
4332: waveform_sig_rx =937;
4333: waveform_sig_rx =1249;
4334: waveform_sig_rx =880;
4335: waveform_sig_rx =1046;
4336: waveform_sig_rx =1214;
4337: waveform_sig_rx =856;
4338: waveform_sig_rx =1035;
4339: waveform_sig_rx =1248;
4340: waveform_sig_rx =847;
4341: waveform_sig_rx =1005;
4342: waveform_sig_rx =1262;
4343: waveform_sig_rx =822;
4344: waveform_sig_rx =1010;
4345: waveform_sig_rx =1188;
4346: waveform_sig_rx =941;
4347: waveform_sig_rx =867;
4348: waveform_sig_rx =1176;
4349: waveform_sig_rx =982;
4350: waveform_sig_rx =911;
4351: waveform_sig_rx =1012;
4352: waveform_sig_rx =1119;
4353: waveform_sig_rx =904;
4354: waveform_sig_rx =941;
4355: waveform_sig_rx =1146;
4356: waveform_sig_rx =926;
4357: waveform_sig_rx =855;
4358: waveform_sig_rx =1162;
4359: waveform_sig_rx =989;
4360: waveform_sig_rx =794;
4361: waveform_sig_rx =1117;
4362: waveform_sig_rx =986;
4363: waveform_sig_rx =816;
4364: waveform_sig_rx =1009;
4365: waveform_sig_rx =1068;
4366: waveform_sig_rx =837;
4367: waveform_sig_rx =986;
4368: waveform_sig_rx =894;
4369: waveform_sig_rx =950;
4370: waveform_sig_rx =931;
4371: waveform_sig_rx =918;
4372: waveform_sig_rx =946;
4373: waveform_sig_rx =779;
4374: waveform_sig_rx =1131;
4375: waveform_sig_rx =711;
4376: waveform_sig_rx =911;
4377: waveform_sig_rx =1072;
4378: waveform_sig_rx =668;
4379: waveform_sig_rx =923;
4380: waveform_sig_rx =1089;
4381: waveform_sig_rx =633;
4382: waveform_sig_rx =898;
4383: waveform_sig_rx =1070;
4384: waveform_sig_rx =623;
4385: waveform_sig_rx =903;
4386: waveform_sig_rx =952;
4387: waveform_sig_rx =780;
4388: waveform_sig_rx =732;
4389: waveform_sig_rx =981;
4390: waveform_sig_rx =832;
4391: waveform_sig_rx =748;
4392: waveform_sig_rx =824;
4393: waveform_sig_rx =999;
4394: waveform_sig_rx =660;
4395: waveform_sig_rx =773;
4396: waveform_sig_rx =1016;
4397: waveform_sig_rx =665;
4398: waveform_sig_rx =697;
4399: waveform_sig_rx =969;
4400: waveform_sig_rx =738;
4401: waveform_sig_rx =653;
4402: waveform_sig_rx =901;
4403: waveform_sig_rx =807;
4404: waveform_sig_rx =645;
4405: waveform_sig_rx =780;
4406: waveform_sig_rx =911;
4407: waveform_sig_rx =625;
4408: waveform_sig_rx =781;
4409: waveform_sig_rx =706;
4410: waveform_sig_rx =757;
4411: waveform_sig_rx =693;
4412: waveform_sig_rx =750;
4413: waveform_sig_rx =705;
4414: waveform_sig_rx =582;
4415: waveform_sig_rx =957;
4416: waveform_sig_rx =448;
4417: waveform_sig_rx =741;
4418: waveform_sig_rx =873;
4419: waveform_sig_rx =402;
4420: waveform_sig_rx =803;
4421: waveform_sig_rx =819;
4422: waveform_sig_rx =411;
4423: waveform_sig_rx =753;
4424: waveform_sig_rx =780;
4425: waveform_sig_rx =480;
4426: waveform_sig_rx =673;
4427: waveform_sig_rx =732;
4428: waveform_sig_rx =605;
4429: waveform_sig_rx =459;
4430: waveform_sig_rx =792;
4431: waveform_sig_rx =600;
4432: waveform_sig_rx =486;
4433: waveform_sig_rx =642;
4434: waveform_sig_rx =728;
4435: waveform_sig_rx =424;
4436: waveform_sig_rx =587;
4437: waveform_sig_rx =744;
4438: waveform_sig_rx =429;
4439: waveform_sig_rx =506;
4440: waveform_sig_rx =703;
4441: waveform_sig_rx =493;
4442: waveform_sig_rx =430;
4443: waveform_sig_rx =620;
4444: waveform_sig_rx =593;
4445: waveform_sig_rx =398;
4446: waveform_sig_rx =506;
4447: waveform_sig_rx =705;
4448: waveform_sig_rx =317;
4449: waveform_sig_rx =540;
4450: waveform_sig_rx =471;
4451: waveform_sig_rx =465;
4452: waveform_sig_rx =471;
4453: waveform_sig_rx =513;
4454: waveform_sig_rx =404;
4455: waveform_sig_rx =402;
4456: waveform_sig_rx =655;
4457: waveform_sig_rx =170;
4458: waveform_sig_rx =556;
4459: waveform_sig_rx =534;
4460: waveform_sig_rx =187;
4461: waveform_sig_rx =544;
4462: waveform_sig_rx =500;
4463: waveform_sig_rx =213;
4464: waveform_sig_rx =468;
4465: waveform_sig_rx =504;
4466: waveform_sig_rx =238;
4467: waveform_sig_rx =381;
4468: waveform_sig_rx =473;
4469: waveform_sig_rx =320;
4470: waveform_sig_rx =184;
4471: waveform_sig_rx =547;
4472: waveform_sig_rx =311;
4473: waveform_sig_rx =204;
4474: waveform_sig_rx =385;
4475: waveform_sig_rx =432;
4476: waveform_sig_rx =129;
4477: waveform_sig_rx =352;
4478: waveform_sig_rx =412;
4479: waveform_sig_rx =153;
4480: waveform_sig_rx =273;
4481: waveform_sig_rx =376;
4482: waveform_sig_rx =275;
4483: waveform_sig_rx =110;
4484: waveform_sig_rx =336;
4485: waveform_sig_rx =326;
4486: waveform_sig_rx =29;
4487: waveform_sig_rx =283;
4488: waveform_sig_rx =388;
4489: waveform_sig_rx =-3;
4490: waveform_sig_rx =329;
4491: waveform_sig_rx =138;
4492: waveform_sig_rx =210;
4493: waveform_sig_rx =205;
4494: waveform_sig_rx =189;
4495: waveform_sig_rx =118;
4496: waveform_sig_rx =134;
4497: waveform_sig_rx =330;
4498: waveform_sig_rx =-86;
4499: waveform_sig_rx =270;
4500: waveform_sig_rx =191;
4501: waveform_sig_rx =-81;
4502: waveform_sig_rx =234;
4503: waveform_sig_rx =183;
4504: waveform_sig_rx =-78;
4505: waveform_sig_rx =137;
4506: waveform_sig_rx =222;
4507: waveform_sig_rx =-72;
4508: waveform_sig_rx =44;
4509: waveform_sig_rx =225;
4510: waveform_sig_rx =-20;
4511: waveform_sig_rx =-122;
4512: waveform_sig_rx =276;
4513: waveform_sig_rx =-58;
4514: waveform_sig_rx =-60;
4515: waveform_sig_rx =94;
4516: waveform_sig_rx =100;
4517: waveform_sig_rx =-130;
4518: waveform_sig_rx =38;
4519: waveform_sig_rx =124;
4520: waveform_sig_rx =-102;
4521: waveform_sig_rx =-100;
4522: waveform_sig_rx =107;
4523: waveform_sig_rx =-33;
4524: waveform_sig_rx =-216;
4525: waveform_sig_rx =104;
4526: waveform_sig_rx =18;
4527: waveform_sig_rx =-257;
4528: waveform_sig_rx =37;
4529: waveform_sig_rx =35;
4530: waveform_sig_rx =-279;
4531: waveform_sig_rx =43;
4532: waveform_sig_rx =-223;
4533: waveform_sig_rx =-61;
4534: waveform_sig_rx =-131;
4535: waveform_sig_rx =-132;
4536: waveform_sig_rx =-167;
4537: waveform_sig_rx =-176;
4538: waveform_sig_rx =3;
4539: waveform_sig_rx =-375;
4540: waveform_sig_rx =-62;
4541: waveform_sig_rx =-80;
4542: waveform_sig_rx =-380;
4543: waveform_sig_rx =-80;
4544: waveform_sig_rx =-71;
4545: waveform_sig_rx =-391;
4546: waveform_sig_rx =-156;
4547: waveform_sig_rx =-54;
4548: waveform_sig_rx =-409;
4549: waveform_sig_rx =-240;
4550: waveform_sig_rx =-64;
4551: waveform_sig_rx =-375;
4552: waveform_sig_rx =-342;
4553: waveform_sig_rx =-58;
4554: waveform_sig_rx =-384;
4555: waveform_sig_rx =-309;
4556: waveform_sig_rx =-265;
4557: waveform_sig_rx =-183;
4558: waveform_sig_rx =-426;
4559: waveform_sig_rx =-307;
4560: waveform_sig_rx =-158;
4561: waveform_sig_rx =-447;
4562: waveform_sig_rx =-395;
4563: waveform_sig_rx =-146;
4564: waveform_sig_rx =-390;
4565: waveform_sig_rx =-503;
4566: waveform_sig_rx =-180;
4567: waveform_sig_rx =-352;
4568: waveform_sig_rx =-558;
4569: waveform_sig_rx =-254;
4570: waveform_sig_rx =-304;
4571: waveform_sig_rx =-561;
4572: waveform_sig_rx =-271;
4573: waveform_sig_rx =-540;
4574: waveform_sig_rx =-314;
4575: waveform_sig_rx =-469;
4576: waveform_sig_rx =-408;
4577: waveform_sig_rx =-447;
4578: waveform_sig_rx =-513;
4579: waveform_sig_rx =-250;
4580: waveform_sig_rx =-683;
4581: waveform_sig_rx =-380;
4582: waveform_sig_rx =-350;
4583: waveform_sig_rx =-733;
4584: waveform_sig_rx =-345;
4585: waveform_sig_rx =-384;
4586: waveform_sig_rx =-743;
4587: waveform_sig_rx =-400;
4588: waveform_sig_rx =-379;
4589: waveform_sig_rx =-710;
4590: waveform_sig_rx =-460;
4591: waveform_sig_rx =-382;
4592: waveform_sig_rx =-655;
4593: waveform_sig_rx =-609;
4594: waveform_sig_rx =-363;
4595: waveform_sig_rx =-644;
4596: waveform_sig_rx =-605;
4597: waveform_sig_rx =-560;
4598: waveform_sig_rx =-440;
4599: waveform_sig_rx =-743;
4600: waveform_sig_rx =-580;
4601: waveform_sig_rx =-400;
4602: waveform_sig_rx =-769;
4603: waveform_sig_rx =-641;
4604: waveform_sig_rx =-403;
4605: waveform_sig_rx =-727;
4606: waveform_sig_rx =-705;
4607: waveform_sig_rx =-473;
4608: waveform_sig_rx =-673;
4609: waveform_sig_rx =-753;
4610: waveform_sig_rx =-594;
4611: waveform_sig_rx =-557;
4612: waveform_sig_rx =-808;
4613: waveform_sig_rx =-590;
4614: waveform_sig_rx =-754;
4615: waveform_sig_rx =-603;
4616: waveform_sig_rx =-757;
4617: waveform_sig_rx =-606;
4618: waveform_sig_rx =-782;
4619: waveform_sig_rx =-730;
4620: waveform_sig_rx =-516;
4621: waveform_sig_rx =-960;
4622: waveform_sig_rx =-586;
4623: waveform_sig_rx =-635;
4624: waveform_sig_rx =-993;
4625: waveform_sig_rx =-564;
4626: waveform_sig_rx =-650;
4627: waveform_sig_rx =-1006;
4628: waveform_sig_rx =-620;
4629: waveform_sig_rx =-673;
4630: waveform_sig_rx =-989;
4631: waveform_sig_rx =-675;
4632: waveform_sig_rx =-707;
4633: waveform_sig_rx =-889;
4634: waveform_sig_rx =-844;
4635: waveform_sig_rx =-679;
4636: waveform_sig_rx =-839;
4637: waveform_sig_rx =-920;
4638: waveform_sig_rx =-780;
4639: waveform_sig_rx =-669;
4640: waveform_sig_rx =-1064;
4641: waveform_sig_rx =-731;
4642: waveform_sig_rx =-710;
4643: waveform_sig_rx =-1044;
4644: waveform_sig_rx =-829;
4645: waveform_sig_rx =-707;
4646: waveform_sig_rx =-922;
4647: waveform_sig_rx =-961;
4648: waveform_sig_rx =-733;
4649: waveform_sig_rx =-867;
4650: waveform_sig_rx =-1028;
4651: waveform_sig_rx =-806;
4652: waveform_sig_rx =-787;
4653: waveform_sig_rx =-1054;
4654: waveform_sig_rx =-823;
4655: waveform_sig_rx =-974;
4656: waveform_sig_rx =-848;
4657: waveform_sig_rx =-974;
4658: waveform_sig_rx =-827;
4659: waveform_sig_rx =-1041;
4660: waveform_sig_rx =-907;
4661: waveform_sig_rx =-772;
4662: waveform_sig_rx =-1207;
4663: waveform_sig_rx =-788;
4664: waveform_sig_rx =-914;
4665: waveform_sig_rx =-1202;
4666: waveform_sig_rx =-764;
4667: waveform_sig_rx =-926;
4668: waveform_sig_rx =-1190;
4669: waveform_sig_rx =-818;
4670: waveform_sig_rx =-945;
4671: waveform_sig_rx =-1153;
4672: waveform_sig_rx =-926;
4673: waveform_sig_rx =-903;
4674: waveform_sig_rx =-1058;
4675: waveform_sig_rx =-1118;
4676: waveform_sig_rx =-807;
4677: waveform_sig_rx =-1060;
4678: waveform_sig_rx =-1158;
4679: waveform_sig_rx =-871;
4680: waveform_sig_rx =-944;
4681: waveform_sig_rx =-1223;
4682: waveform_sig_rx =-891;
4683: waveform_sig_rx =-961;
4684: waveform_sig_rx =-1135;
4685: waveform_sig_rx =-1055;
4686: waveform_sig_rx =-901;
4687: waveform_sig_rx =-1080;
4688: waveform_sig_rx =-1164;
4689: waveform_sig_rx =-857;
4690: waveform_sig_rx =-1069;
4691: waveform_sig_rx =-1185;
4692: waveform_sig_rx =-947;
4693: waveform_sig_rx =-977;
4694: waveform_sig_rx =-1190;
4695: waveform_sig_rx =-997;
4696: waveform_sig_rx =-1107;
4697: waveform_sig_rx =-1026;
4698: waveform_sig_rx =-1108;
4699: waveform_sig_rx =-973;
4700: waveform_sig_rx =-1230;
4701: waveform_sig_rx =-986;
4702: waveform_sig_rx =-993;
4703: waveform_sig_rx =-1331;
4704: waveform_sig_rx =-871;
4705: waveform_sig_rx =-1136;
4706: waveform_sig_rx =-1225;
4707: waveform_sig_rx =-941;
4708: waveform_sig_rx =-1074;
4709: waveform_sig_rx =-1261;
4710: waveform_sig_rx =-1031;
4711: waveform_sig_rx =-1001;
4712: waveform_sig_rx =-1294;
4713: waveform_sig_rx =-1061;
4714: waveform_sig_rx =-960;
4715: waveform_sig_rx =-1260;
4716: waveform_sig_rx =-1192;
4717: waveform_sig_rx =-930;
4718: waveform_sig_rx =-1215;
4719: waveform_sig_rx =-1202;
4720: waveform_sig_rx =-1026;
4721: waveform_sig_rx =-1072;
4722: waveform_sig_rx =-1302;
4723: waveform_sig_rx =-1034;
4724: waveform_sig_rx =-1071;
4725: waveform_sig_rx =-1263;
4726: waveform_sig_rx =-1138;
4727: waveform_sig_rx =-1003;
4728: waveform_sig_rx =-1208;
4729: waveform_sig_rx =-1266;
4730: waveform_sig_rx =-984;
4731: waveform_sig_rx =-1162;
4732: waveform_sig_rx =-1313;
4733: waveform_sig_rx =-1012;
4734: waveform_sig_rx =-1092;
4735: waveform_sig_rx =-1323;
4736: waveform_sig_rx =-1012;
4737: waveform_sig_rx =-1262;
4738: waveform_sig_rx =-1094;
4739: waveform_sig_rx =-1162;
4740: waveform_sig_rx =-1119;
4741: waveform_sig_rx =-1269;
4742: waveform_sig_rx =-1072;
4743: waveform_sig_rx =-1129;
4744: waveform_sig_rx =-1323;
4745: waveform_sig_rx =-1019;
4746: waveform_sig_rx =-1173;
4747: waveform_sig_rx =-1290;
4748: waveform_sig_rx =-1043;
4749: waveform_sig_rx =-1075;
4750: waveform_sig_rx =-1403;
4751: waveform_sig_rx =-1011;
4752: waveform_sig_rx =-1076;
4753: waveform_sig_rx =-1396;
4754: waveform_sig_rx =-1049;
4755: waveform_sig_rx =-1066;
4756: waveform_sig_rx =-1295;
4757: waveform_sig_rx =-1179;
4758: waveform_sig_rx =-984;
4759: waveform_sig_rx =-1242;
4760: waveform_sig_rx =-1236;
4761: waveform_sig_rx =-1051;
4762: waveform_sig_rx =-1131;
4763: waveform_sig_rx =-1302;
4764: waveform_sig_rx =-1052;
4765: waveform_sig_rx =-1122;
4766: waveform_sig_rx =-1265;
4767: waveform_sig_rx =-1205;
4768: waveform_sig_rx =-987;
4769: waveform_sig_rx =-1244;
4770: waveform_sig_rx =-1316;
4771: waveform_sig_rx =-903;
4772: waveform_sig_rx =-1258;
4773: waveform_sig_rx =-1284;
4774: waveform_sig_rx =-973;
4775: waveform_sig_rx =-1174;
4776: waveform_sig_rx =-1235;
4777: waveform_sig_rx =-1056;
4778: waveform_sig_rx =-1274;
4779: waveform_sig_rx =-1008;
4780: waveform_sig_rx =-1233;
4781: waveform_sig_rx =-1064;
4782: waveform_sig_rx =-1246;
4783: waveform_sig_rx =-1104;
4784: waveform_sig_rx =-1048;
4785: waveform_sig_rx =-1326;
4786: waveform_sig_rx =-980;
4787: waveform_sig_rx =-1106;
4788: waveform_sig_rx =-1334;
4789: waveform_sig_rx =-945;
4790: waveform_sig_rx =-1075;
4791: waveform_sig_rx =-1352;
4792: waveform_sig_rx =-935;
4793: waveform_sig_rx =-1062;
4794: waveform_sig_rx =-1318;
4795: waveform_sig_rx =-980;
4796: waveform_sig_rx =-1028;
4797: waveform_sig_rx =-1268;
4798: waveform_sig_rx =-1114;
4799: waveform_sig_rx =-960;
4800: waveform_sig_rx =-1209;
4801: waveform_sig_rx =-1152;
4802: waveform_sig_rx =-1018;
4803: waveform_sig_rx =-1062;
4804: waveform_sig_rx =-1225;
4805: waveform_sig_rx =-1043;
4806: waveform_sig_rx =-975;
4807: waveform_sig_rx =-1246;
4808: waveform_sig_rx =-1117;
4809: waveform_sig_rx =-851;
4810: waveform_sig_rx =-1258;
4811: waveform_sig_rx =-1136;
4812: waveform_sig_rx =-866;
4813: waveform_sig_rx =-1200;
4814: waveform_sig_rx =-1119;
4815: waveform_sig_rx =-961;
4816: waveform_sig_rx =-1045;
4817: waveform_sig_rx =-1133;
4818: waveform_sig_rx =-1004;
4819: waveform_sig_rx =-1108;
4820: waveform_sig_rx =-983;
4821: waveform_sig_rx =-1131;
4822: waveform_sig_rx =-927;
4823: waveform_sig_rx =-1207;
4824: waveform_sig_rx =-956;
4825: waveform_sig_rx =-988;
4826: waveform_sig_rx =-1249;
4827: waveform_sig_rx =-852;
4828: waveform_sig_rx =-1053;
4829: waveform_sig_rx =-1216;
4830: waveform_sig_rx =-829;
4831: waveform_sig_rx =-992;
4832: waveform_sig_rx =-1268;
4833: waveform_sig_rx =-786;
4834: waveform_sig_rx =-998;
4835: waveform_sig_rx =-1212;
4836: waveform_sig_rx =-817;
4837: waveform_sig_rx =-964;
4838: waveform_sig_rx =-1114;
4839: waveform_sig_rx =-960;
4840: waveform_sig_rx =-874;
4841: waveform_sig_rx =-1040;
4842: waveform_sig_rx =-1056;
4843: waveform_sig_rx =-864;
4844: waveform_sig_rx =-888;
4845: waveform_sig_rx =-1178;
4846: waveform_sig_rx =-796;
4847: waveform_sig_rx =-868;
4848: waveform_sig_rx =-1144;
4849: waveform_sig_rx =-894;
4850: waveform_sig_rx =-788;
4851: waveform_sig_rx =-1085;
4852: waveform_sig_rx =-936;
4853: waveform_sig_rx =-753;
4854: waveform_sig_rx =-997;
4855: waveform_sig_rx =-997;
4856: waveform_sig_rx =-812;
4857: waveform_sig_rx =-859;
4858: waveform_sig_rx =-1015;
4859: waveform_sig_rx =-818;
4860: waveform_sig_rx =-931;
4861: waveform_sig_rx =-825;
4862: waveform_sig_rx =-943;
4863: waveform_sig_rx =-739;
4864: waveform_sig_rx =-1061;
4865: waveform_sig_rx =-720;
4866: waveform_sig_rx =-815;
4867: waveform_sig_rx =-1061;
4868: waveform_sig_rx =-640;
4869: waveform_sig_rx =-919;
4870: waveform_sig_rx =-1006;
4871: waveform_sig_rx =-622;
4872: waveform_sig_rx =-868;
4873: waveform_sig_rx =-1017;
4874: waveform_sig_rx =-596;
4875: waveform_sig_rx =-857;
4876: waveform_sig_rx =-961;
4877: waveform_sig_rx =-692;
4878: waveform_sig_rx =-787;
4879: waveform_sig_rx =-924;
4880: waveform_sig_rx =-824;
4881: waveform_sig_rx =-651;
4882: waveform_sig_rx =-847;
4883: waveform_sig_rx =-881;
4884: waveform_sig_rx =-627;
4885: waveform_sig_rx =-745;
4886: waveform_sig_rx =-972;
4887: waveform_sig_rx =-573;
4888: waveform_sig_rx =-736;
4889: waveform_sig_rx =-907;
4890: waveform_sig_rx =-679;
4891: waveform_sig_rx =-643;
4892: waveform_sig_rx =-855;
4893: waveform_sig_rx =-754;
4894: waveform_sig_rx =-588;
4895: waveform_sig_rx =-751;
4896: waveform_sig_rx =-836;
4897: waveform_sig_rx =-566;
4898: waveform_sig_rx =-663;
4899: waveform_sig_rx =-832;
4900: waveform_sig_rx =-561;
4901: waveform_sig_rx =-759;
4902: waveform_sig_rx =-612;
4903: waveform_sig_rx =-708;
4904: waveform_sig_rx =-557;
4905: waveform_sig_rx =-836;
4906: waveform_sig_rx =-484;
4907: waveform_sig_rx =-649;
4908: waveform_sig_rx =-823;
4909: waveform_sig_rx =-383;
4910: waveform_sig_rx =-738;
4911: waveform_sig_rx =-737;
4912: waveform_sig_rx =-391;
4913: waveform_sig_rx =-683;
4914: waveform_sig_rx =-734;
4915: waveform_sig_rx =-403;
4916: waveform_sig_rx =-628;
4917: waveform_sig_rx =-679;
4918: waveform_sig_rx =-474;
4919: waveform_sig_rx =-486;
4920: waveform_sig_rx =-704;
4921: waveform_sig_rx =-559;
4922: waveform_sig_rx =-376;
4923: waveform_sig_rx =-667;
4924: waveform_sig_rx =-612;
4925: waveform_sig_rx =-377;
4926: waveform_sig_rx =-532;
4927: waveform_sig_rx =-675;
4928: waveform_sig_rx =-341;
4929: waveform_sig_rx =-498;
4930: waveform_sig_rx =-605;
4931: waveform_sig_rx =-448;
4932: waveform_sig_rx =-380;
4933: waveform_sig_rx =-570;
4934: waveform_sig_rx =-550;
4935: waveform_sig_rx =-307;
4936: waveform_sig_rx =-520;
4937: waveform_sig_rx =-602;
4938: waveform_sig_rx =-249;
4939: waveform_sig_rx =-444;
4940: waveform_sig_rx =-551;
4941: waveform_sig_rx =-289;
4942: waveform_sig_rx =-550;
4943: waveform_sig_rx =-294;
4944: waveform_sig_rx =-456;
4945: waveform_sig_rx =-311;
4946: waveform_sig_rx =-534;
4947: waveform_sig_rx =-202;
4948: waveform_sig_rx =-400;
4949: waveform_sig_rx =-521;
4950: waveform_sig_rx =-132;
4951: waveform_sig_rx =-462;
4952: waveform_sig_rx =-447;
4953: waveform_sig_rx =-126;
4954: waveform_sig_rx =-402;
4955: waveform_sig_rx =-453;
4956: waveform_sig_rx =-159;
4957: waveform_sig_rx =-309;
4958: waveform_sig_rx =-415;
4959: waveform_sig_rx =-234;
4960: waveform_sig_rx =-173;
4961: waveform_sig_rx =-511;
4962: waveform_sig_rx =-214;
4963: waveform_sig_rx =-111;
4964: waveform_sig_rx =-422;
4965: waveform_sig_rx =-237;
4966: waveform_sig_rx =-153;
4967: waveform_sig_rx =-251;
4968: waveform_sig_rx =-348;
4969: waveform_sig_rx =-109;
4970: waveform_sig_rx =-162;
4971: waveform_sig_rx =-361;
4972: waveform_sig_rx =-141;
4973: waveform_sig_rx =-53;
4974: waveform_sig_rx =-341;
4975: waveform_sig_rx =-206;
4976: waveform_sig_rx =1;
4977: waveform_sig_rx =-257;
4978: waveform_sig_rx =-282;
4979: waveform_sig_rx =25;
4980: waveform_sig_rx =-204;
4981: waveform_sig_rx =-240;
4982: waveform_sig_rx =-10;
4983: waveform_sig_rx =-252;
4984: waveform_sig_rx =9;
4985: waveform_sig_rx =-174;
4986: waveform_sig_rx =-29;
4987: waveform_sig_rx =-246;
4988: waveform_sig_rx =45;
4989: waveform_sig_rx =-128;
4990: waveform_sig_rx =-189;
4991: waveform_sig_rx =108;
4992: waveform_sig_rx =-149;
4993: waveform_sig_rx =-166;
4994: waveform_sig_rx =142;
4995: waveform_sig_rx =-75;
4996: waveform_sig_rx =-204;
4997: waveform_sig_rx =177;
4998: waveform_sig_rx =-38;
4999: waveform_sig_rx =-185;
5000: waveform_sig_rx =128;
5001: waveform_sig_rx =55;
5002: waveform_sig_rx =-210;
5003: waveform_sig_rx =134;
5004: waveform_sig_rx =107;
5005: waveform_sig_rx =-81;
5006: waveform_sig_rx =26;
5007: waveform_sig_rx =129;
5008: waveform_sig_rx =88;
5009: waveform_sig_rx =-102;
5010: waveform_sig_rx =203;
5011: waveform_sig_rx =128;
5012: waveform_sig_rx =-87;
5013: waveform_sig_rx =167;
5014: waveform_sig_rx =215;
5015: waveform_sig_rx =-58;
5016: waveform_sig_rx =88;
5017: waveform_sig_rx =300;
5018: waveform_sig_rx =-20;
5019: waveform_sig_rx =44;
5020: waveform_sig_rx =322;
5021: waveform_sig_rx =64;
5022: waveform_sig_rx =120;
5023: waveform_sig_rx =226;
5024: waveform_sig_rx =63;
5025: waveform_sig_rx =304;
5026: waveform_sig_rx =68;
5027: waveform_sig_rx =300;
5028: waveform_sig_rx =31;
5029: waveform_sig_rx =341;
5030: waveform_sig_rx =216;
5031: waveform_sig_rx =51;
5032: waveform_sig_rx =439;
5033: waveform_sig_rx =161;
5034: waveform_sig_rx =97;
5035: waveform_sig_rx =520;
5036: waveform_sig_rx =152;
5037: waveform_sig_rx =94;
5038: waveform_sig_rx =512;
5039: waveform_sig_rx =187;
5040: waveform_sig_rx =161;
5041: waveform_sig_rx =426;
5042: waveform_sig_rx =332;
5043: waveform_sig_rx =121;
5044: waveform_sig_rx =408;
5045: waveform_sig_rx =376;
5046: waveform_sig_rx =236;
5047: waveform_sig_rx =294;
5048: waveform_sig_rx =427;
5049: waveform_sig_rx =352;
5050: waveform_sig_rx =158;
5051: waveform_sig_rx =520;
5052: waveform_sig_rx =391;
5053: waveform_sig_rx =174;
5054: waveform_sig_rx =498;
5055: waveform_sig_rx =480;
5056: waveform_sig_rx =208;
5057: waveform_sig_rx =435;
5058: waveform_sig_rx =542;
5059: waveform_sig_rx =288;
5060: waveform_sig_rx =369;
5061: waveform_sig_rx =555;
5062: waveform_sig_rx =358;
5063: waveform_sig_rx =387;
5064: waveform_sig_rx =451;
5065: waveform_sig_rx =390;
5066: waveform_sig_rx =524;
5067: waveform_sig_rx =371;
5068: waveform_sig_rx =602;
5069: waveform_sig_rx =265;
5070: waveform_sig_rx =677;
5071: waveform_sig_rx =441;
5072: waveform_sig_rx =309;
5073: waveform_sig_rx =752;
5074: waveform_sig_rx =357;
5075: waveform_sig_rx =410;
5076: waveform_sig_rx =785;
5077: waveform_sig_rx =391;
5078: waveform_sig_rx =411;
5079: waveform_sig_rx =768;
5080: waveform_sig_rx =451;
5081: waveform_sig_rx =444;
5082: waveform_sig_rx =690;
5083: waveform_sig_rx =588;
5084: waveform_sig_rx =392;
5085: waveform_sig_rx =670;
5086: waveform_sig_rx =643;
5087: waveform_sig_rx =509;
5088: waveform_sig_rx =530;
5089: waveform_sig_rx =742;
5090: waveform_sig_rx =602;
5091: waveform_sig_rx =408;
5092: waveform_sig_rx =844;
5093: waveform_sig_rx =587;
5094: waveform_sig_rx =452;
5095: waveform_sig_rx =804;
5096: waveform_sig_rx =667;
5097: waveform_sig_rx =519;
5098: waveform_sig_rx =681;
5099: waveform_sig_rx =753;
5100: waveform_sig_rx =598;
5101: waveform_sig_rx =571;
5102: waveform_sig_rx =851;
5103: waveform_sig_rx =638;
5104: waveform_sig_rx =598;
5105: waveform_sig_rx =758;
5106: waveform_sig_rx =637;
5107: waveform_sig_rx =760;
5108: waveform_sig_rx =666;
5109: waveform_sig_rx =799;
5110: waveform_sig_rx =505;
5111: waveform_sig_rx =954;
5112: waveform_sig_rx =622;
5113: waveform_sig_rx =584;
5114: waveform_sig_rx =1022;
5115: waveform_sig_rx =550;
5116: waveform_sig_rx =671;
5117: waveform_sig_rx =1012;
5118: waveform_sig_rx =576;
5119: waveform_sig_rx =716;
5120: waveform_sig_rx =978;
5121: waveform_sig_rx =648;
5122: waveform_sig_rx =736;
5123: waveform_sig_rx =866;
5124: waveform_sig_rx =845;
5125: waveform_sig_rx =644;
5126: waveform_sig_rx =869;
5127: waveform_sig_rx =925;
5128: waveform_sig_rx =696;
5129: waveform_sig_rx =769;
5130: waveform_sig_rx =993;
5131: waveform_sig_rx =725;
5132: waveform_sig_rx =717;
5133: waveform_sig_rx =1055;
5134: waveform_sig_rx =784;
5135: waveform_sig_rx =733;
5136: waveform_sig_rx =959;
5137: waveform_sig_rx =910;
5138: waveform_sig_rx =739;
5139: waveform_sig_rx =877;
5140: waveform_sig_rx =1006;
5141: waveform_sig_rx =793;
5142: waveform_sig_rx =792;
5143: waveform_sig_rx =1084;
5144: waveform_sig_rx =820;
5145: waveform_sig_rx =819;
5146: waveform_sig_rx =987;
5147: waveform_sig_rx =846;
5148: waveform_sig_rx =952;
5149: waveform_sig_rx =917;
5150: waveform_sig_rx =966;
5151: waveform_sig_rx =748;
5152: waveform_sig_rx =1199;
5153: waveform_sig_rx =766;
5154: waveform_sig_rx =886;
5155: waveform_sig_rx =1168;
5156: waveform_sig_rx =734;
5157: waveform_sig_rx =959;
5158: waveform_sig_rx =1136;
5159: waveform_sig_rx =826;
5160: waveform_sig_rx =904;
5161: waveform_sig_rx =1119;
5162: waveform_sig_rx =893;
5163: waveform_sig_rx =894;
5164: waveform_sig_rx =1080;
5165: waveform_sig_rx =1051;
5166: waveform_sig_rx =780;
5167: waveform_sig_rx =1104;
5168: waveform_sig_rx =1093;
5169: waveform_sig_rx =852;
5170: waveform_sig_rx =1005;
5171: waveform_sig_rx =1174;
5172: waveform_sig_rx =904;
5173: waveform_sig_rx =912;
5174: waveform_sig_rx =1187;
5175: waveform_sig_rx =964;
5176: waveform_sig_rx =924;
5177: waveform_sig_rx =1122;
5178: waveform_sig_rx =1103;
5179: waveform_sig_rx =895;
5180: waveform_sig_rx =1028;
5181: waveform_sig_rx =1193;
5182: waveform_sig_rx =905;
5183: waveform_sig_rx =962;
5184: waveform_sig_rx =1285;
5185: waveform_sig_rx =931;
5186: waveform_sig_rx =1002;
5187: waveform_sig_rx =1159;
5188: waveform_sig_rx =937;
5189: waveform_sig_rx =1152;
5190: waveform_sig_rx =1057;
5191: waveform_sig_rx =1056;
5192: waveform_sig_rx =948;
5193: waveform_sig_rx =1262;
5194: waveform_sig_rx =891;
5195: waveform_sig_rx =1077;
5196: waveform_sig_rx =1224;
5197: waveform_sig_rx =946;
5198: waveform_sig_rx =1071;
5199: waveform_sig_rx =1251;
5200: waveform_sig_rx =993;
5201: waveform_sig_rx =964;
5202: waveform_sig_rx =1325;
5203: waveform_sig_rx =970;
5204: waveform_sig_rx =1004;
5205: waveform_sig_rx =1260;
5206: waveform_sig_rx =1099;
5207: waveform_sig_rx =923;
5208: waveform_sig_rx =1230;
5209: waveform_sig_rx =1167;
5210: waveform_sig_rx =967;
5211: waveform_sig_rx =1108;
5212: waveform_sig_rx =1276;
5213: waveform_sig_rx =982;
5214: waveform_sig_rx =1080;
5215: waveform_sig_rx =1250;
5216: waveform_sig_rx =1075;
5217: waveform_sig_rx =1043;
5218: waveform_sig_rx =1180;
5219: waveform_sig_rx =1278;
5220: waveform_sig_rx =898;
5221: waveform_sig_rx =1178;
5222: waveform_sig_rx =1316;
5223: waveform_sig_rx =896;
5224: waveform_sig_rx =1163;
5225: waveform_sig_rx =1306;
5226: waveform_sig_rx =964;
5227: waveform_sig_rx =1199;
5228: waveform_sig_rx =1121;
5229: waveform_sig_rx =1093;
5230: waveform_sig_rx =1218;
5231: waveform_sig_rx =1080;
5232: waveform_sig_rx =1210;
5233: waveform_sig_rx =1016;
5234: waveform_sig_rx =1318;
5235: waveform_sig_rx =1018;
5236: waveform_sig_rx =1107;
5237: waveform_sig_rx =1310;
5238: waveform_sig_rx =1021;
5239: waveform_sig_rx =1109;
5240: waveform_sig_rx =1354;
5241: waveform_sig_rx =1017;
5242: waveform_sig_rx =1044;
5243: waveform_sig_rx =1415;
5244: waveform_sig_rx =995;
5245: waveform_sig_rx =1049;
5246: waveform_sig_rx =1329;
5247: waveform_sig_rx =1113;
5248: waveform_sig_rx =980;
5249: waveform_sig_rx =1304;
5250: waveform_sig_rx =1150;
5251: waveform_sig_rx =1042;
5252: waveform_sig_rx =1164;
5253: waveform_sig_rx =1252;
5254: waveform_sig_rx =1057;
5255: waveform_sig_rx =1071;
5256: waveform_sig_rx =1271;
5257: waveform_sig_rx =1150;
5258: waveform_sig_rx =980;
5259: waveform_sig_rx =1273;
5260: waveform_sig_rx =1253;
5261: waveform_sig_rx =901;
5262: waveform_sig_rx =1297;
5263: waveform_sig_rx =1248;
5264: waveform_sig_rx =972;
5265: waveform_sig_rx =1222;
5266: waveform_sig_rx =1255;
5267: waveform_sig_rx =1058;
5268: waveform_sig_rx =1161;
5269: waveform_sig_rx =1123;
5270: waveform_sig_rx =1166;
5271: waveform_sig_rx =1188;
5272: waveform_sig_rx =1123;
5273: waveform_sig_rx =1205;
5274: waveform_sig_rx =985;
5275: waveform_sig_rx =1354;
5276: waveform_sig_rx =986;
5277: waveform_sig_rx =1103;
5278: waveform_sig_rx =1328;
5279: waveform_sig_rx =985;
5280: waveform_sig_rx =1093;
5281: waveform_sig_rx =1363;
5282: waveform_sig_rx =978;
5283: waveform_sig_rx =1041;
5284: waveform_sig_rx =1425;
5285: waveform_sig_rx =921;
5286: waveform_sig_rx =1117;
5287: waveform_sig_rx =1307;
5288: waveform_sig_rx =1040;
5289: waveform_sig_rx =1016;
5290: waveform_sig_rx =1244;
5291: waveform_sig_rx =1132;
5292: waveform_sig_rx =1045;
5293: waveform_sig_rx =1087;
5294: waveform_sig_rx =1288;
5295: waveform_sig_rx =1019;
5296: waveform_sig_rx =1022;
5297: waveform_sig_rx =1316;
5298: waveform_sig_rx =1028;
5299: waveform_sig_rx =971;
5300: waveform_sig_rx =1282;
5301: waveform_sig_rx =1118;
5302: waveform_sig_rx =928;
5303: waveform_sig_rx =1238;
5304: waveform_sig_rx =1149;
5305: waveform_sig_rx =970;
5306: waveform_sig_rx =1098;
5307: waveform_sig_rx =1231;
5308: waveform_sig_rx =1004;
5309: waveform_sig_rx =1076;
5310: waveform_sig_rx =1085;
5311: waveform_sig_rx =1082;
5312: waveform_sig_rx =1079;
5313: waveform_sig_rx =1088;
5314: waveform_sig_rx =1117;
5315: waveform_sig_rx =908;
5316: waveform_sig_rx =1305;
5317: waveform_sig_rx =883;
5318: waveform_sig_rx =1029;
5319: waveform_sig_rx =1277;
5320: waveform_sig_rx =843;
5321: waveform_sig_rx =1060;
5322: waveform_sig_rx =1301;
5323: waveform_sig_rx =813;
5324: waveform_sig_rx =1051;
5325: waveform_sig_rx =1261;
5326: waveform_sig_rx =820;
5327: waveform_sig_rx =1072;
5328: waveform_sig_rx =1140;
5329: waveform_sig_rx =990;
5330: waveform_sig_rx =899;
5331: waveform_sig_rx =1103;
5332: waveform_sig_rx =1065;
5333: waveform_sig_rx =904;
5334: waveform_sig_rx =977;
5335: waveform_sig_rx =1195;
5336: waveform_sig_rx =832;
5337: waveform_sig_rx =954;
5338: waveform_sig_rx =1188;
5339: waveform_sig_rx =857;
5340: waveform_sig_rx =918;
5341: waveform_sig_rx =1132;
5342: waveform_sig_rx =967;
5343: waveform_sig_rx =831;
5344: waveform_sig_rx =1052;
5345: waveform_sig_rx =1035;
5346: waveform_sig_rx =849;
5347: waveform_sig_rx =940;
5348: waveform_sig_rx =1107;
5349: waveform_sig_rx =834;
5350: waveform_sig_rx =929;
5351: waveform_sig_rx =977;
5352: waveform_sig_rx =915;
5353: waveform_sig_rx =940;
5354: waveform_sig_rx =976;
5355: waveform_sig_rx =897;
5356: waveform_sig_rx =820;
5357: waveform_sig_rx =1164;
5358: waveform_sig_rx =656;
5359: waveform_sig_rx =948;
5360: waveform_sig_rx =1072;
5361: waveform_sig_rx =675;
5362: waveform_sig_rx =960;
5363: waveform_sig_rx =1055;
5364: waveform_sig_rx =673;
5365: waveform_sig_rx =910;
5366: waveform_sig_rx =1034;
5367: waveform_sig_rx =699;
5368: waveform_sig_rx =884;
5369: waveform_sig_rx =930;
5370: waveform_sig_rx =865;
5371: waveform_sig_rx =681;
5372: waveform_sig_rx =968;
5373: waveform_sig_rx =906;
5374: waveform_sig_rx =678;
5375: waveform_sig_rx =879;
5376: waveform_sig_rx =989;
5377: waveform_sig_rx =630;
5378: waveform_sig_rx =861;
5379: waveform_sig_rx =953;
5380: waveform_sig_rx =711;
5381: waveform_sig_rx =761;
5382: waveform_sig_rx =893;
5383: waveform_sig_rx =826;
5384: waveform_sig_rx =629;
5385: waveform_sig_rx =842;
5386: waveform_sig_rx =879;
5387: waveform_sig_rx =609;
5388: waveform_sig_rx =772;
5389: waveform_sig_rx =951;
5390: waveform_sig_rx =583;
5391: waveform_sig_rx =788;
5392: waveform_sig_rx =762;
5393: waveform_sig_rx =691;
5394: waveform_sig_rx =771;
5395: waveform_sig_rx =739;
5396: waveform_sig_rx =668;
5397: waveform_sig_rx =640;
5398: waveform_sig_rx =893;
5399: waveform_sig_rx =452;
5400: waveform_sig_rx =780;
5401: waveform_sig_rx =779;
5402: waveform_sig_rx =490;
5403: waveform_sig_rx =760;
5404: waveform_sig_rx =781;
5405: waveform_sig_rx =507;
5406: waveform_sig_rx =662;
5407: waveform_sig_rx =795;
5408: waveform_sig_rx =514;
5409: waveform_sig_rx =595;
5410: waveform_sig_rx =770;
5411: waveform_sig_rx =610;
5412: waveform_sig_rx =413;
5413: waveform_sig_rx =813;
5414: waveform_sig_rx =605;
5415: waveform_sig_rx =461;
5416: waveform_sig_rx =666;
5417: waveform_sig_rx =685;
5418: waveform_sig_rx =443;
5419: waveform_sig_rx =589;
5420: waveform_sig_rx =696;
5421: waveform_sig_rx =487;
5422: waveform_sig_rx =473;
5423: waveform_sig_rx =674;
5424: waveform_sig_rx =584;
5425: waveform_sig_rx =357;
5426: waveform_sig_rx =647;
5427: waveform_sig_rx =626;
5428: waveform_sig_rx =347;
5429: waveform_sig_rx =563;
5430: waveform_sig_rx =680;
5431: waveform_sig_rx =297;
5432: waveform_sig_rx =582;
5433: waveform_sig_rx =456;
5434: waveform_sig_rx =451;
5435: waveform_sig_rx =541;
5436: waveform_sig_rx =451;
5437: waveform_sig_rx =445;
5438: waveform_sig_rx =399;
5439: waveform_sig_rx =600;
5440: waveform_sig_rx =237;
5441: waveform_sig_rx =503;
5442: waveform_sig_rx =514;
5443: waveform_sig_rx =270;
5444: waveform_sig_rx =439;
5445: waveform_sig_rx =537;
5446: waveform_sig_rx =227;
5447: waveform_sig_rx =364;
5448: waveform_sig_rx =585;
5449: waveform_sig_rx =191;
5450: waveform_sig_rx =338;
5451: waveform_sig_rx =559;
5452: waveform_sig_rx =261;
5453: waveform_sig_rx =197;
5454: waveform_sig_rx =549;
5455: waveform_sig_rx =251;
5456: waveform_sig_rx =269;
5457: waveform_sig_rx =359;
5458: waveform_sig_rx =422;
5459: waveform_sig_rx =169;
5460: waveform_sig_rx =249;
5461: waveform_sig_rx =436;
5462: waveform_sig_rx =173;
5463: waveform_sig_rx =178;
5464: waveform_sig_rx =421;
5465: waveform_sig_rx =260;
5466: waveform_sig_rx =78;
5467: waveform_sig_rx =357;
5468: waveform_sig_rx =326;
5469: waveform_sig_rx =1;
5470: waveform_sig_rx =305;
5471: waveform_sig_rx =363;
5472: waveform_sig_rx =-2;
5473: waveform_sig_rx =360;
5474: waveform_sig_rx =77;
5475: waveform_sig_rx =232;
5476: waveform_sig_rx =220;
5477: waveform_sig_rx =117;
5478: waveform_sig_rx =213;
5479: waveform_sig_rx =49;
5480: waveform_sig_rx =332;
5481: waveform_sig_rx =-16;
5482: waveform_sig_rx =143;
5483: waveform_sig_rx =297;
5484: waveform_sig_rx =-102;
5485: waveform_sig_rx =170;
5486: waveform_sig_rx =312;
5487: waveform_sig_rx =-168;
5488: waveform_sig_rx =149;
5489: waveform_sig_rx =261;
5490: waveform_sig_rx =-123;
5491: waveform_sig_rx =93;
5492: waveform_sig_rx =197;
5493: waveform_sig_rx =-34;
5494: waveform_sig_rx =-81;
5495: waveform_sig_rx =240;
5496: waveform_sig_rx =-48;
5497: waveform_sig_rx =-31;
5498: waveform_sig_rx =37;
5499: waveform_sig_rx =124;
5500: waveform_sig_rx =-125;
5501: waveform_sig_rx =-52;
5502: waveform_sig_rx =171;
5503: waveform_sig_rx =-150;
5504: waveform_sig_rx =-134;
5505: waveform_sig_rx =173;
5506: waveform_sig_rx =-100;
5507: waveform_sig_rx =-219;
5508: waveform_sig_rx =116;
5509: waveform_sig_rx =-59;
5510: waveform_sig_rx =-221;
5511: waveform_sig_rx =0;
5512: waveform_sig_rx =-1;
5513: waveform_sig_rx =-244;
5514: waveform_sig_rx =-33;
5515: waveform_sig_rx =-194;
5516: waveform_sig_rx =-23;
5517: waveform_sig_rx =-166;
5518: waveform_sig_rx =-103;
5519: waveform_sig_rx =-142;
5520: waveform_sig_rx =-275;
5521: waveform_sig_rx =87;
5522: waveform_sig_rx =-420;
5523: waveform_sig_rx =-116;
5524: waveform_sig_rx =-2;
5525: waveform_sig_rx =-461;
5526: waveform_sig_rx =-54;
5527: waveform_sig_rx =-77;
5528: waveform_sig_rx =-463;
5529: waveform_sig_rx =-114;
5530: waveform_sig_rx =-101;
5531: waveform_sig_rx =-408;
5532: waveform_sig_rx =-211;
5533: waveform_sig_rx =-129;
5534: waveform_sig_rx =-374;
5535: waveform_sig_rx =-380;
5536: waveform_sig_rx =-97;
5537: waveform_sig_rx =-348;
5538: waveform_sig_rx =-325;
5539: waveform_sig_rx =-313;
5540: waveform_sig_rx =-141;
5541: waveform_sig_rx =-462;
5542: waveform_sig_rx =-354;
5543: waveform_sig_rx =-100;
5544: waveform_sig_rx =-523;
5545: waveform_sig_rx =-376;
5546: waveform_sig_rx =-144;
5547: waveform_sig_rx =-464;
5548: waveform_sig_rx =-428;
5549: waveform_sig_rx =-265;
5550: waveform_sig_rx =-358;
5551: waveform_sig_rx =-499;
5552: waveform_sig_rx =-376;
5553: waveform_sig_rx =-232;
5554: waveform_sig_rx =-568;
5555: waveform_sig_rx =-355;
5556: waveform_sig_rx =-441;
5557: waveform_sig_rx =-382;
5558: waveform_sig_rx =-457;
5559: waveform_sig_rx =-338;
5560: waveform_sig_rx =-500;
5561: waveform_sig_rx =-501;
5562: waveform_sig_rx =-234;
5563: waveform_sig_rx =-735;
5564: waveform_sig_rx =-340;
5565: waveform_sig_rx =-354;
5566: waveform_sig_rx =-741;
5567: waveform_sig_rx =-327;
5568: waveform_sig_rx =-388;
5569: waveform_sig_rx =-758;
5570: waveform_sig_rx =-389;
5571: waveform_sig_rx =-424;
5572: waveform_sig_rx =-716;
5573: waveform_sig_rx =-457;
5574: waveform_sig_rx =-436;
5575: waveform_sig_rx =-603;
5576: waveform_sig_rx =-678;
5577: waveform_sig_rx =-409;
5578: waveform_sig_rx =-564;
5579: waveform_sig_rx =-702;
5580: waveform_sig_rx =-531;
5581: waveform_sig_rx =-419;
5582: waveform_sig_rx =-821;
5583: waveform_sig_rx =-507;
5584: waveform_sig_rx =-441;
5585: waveform_sig_rx =-774;
5586: waveform_sig_rx =-589;
5587: waveform_sig_rx =-499;
5588: waveform_sig_rx =-659;
5589: waveform_sig_rx =-732;
5590: waveform_sig_rx =-523;
5591: waveform_sig_rx =-571;
5592: waveform_sig_rx =-815;
5593: waveform_sig_rx =-594;
5594: waveform_sig_rx =-526;
5595: waveform_sig_rx =-852;
5596: waveform_sig_rx =-572;
5597: waveform_sig_rx =-732;
5598: waveform_sig_rx =-659;
5599: waveform_sig_rx =-732;
5600: waveform_sig_rx =-641;
5601: waveform_sig_rx =-815;
5602: waveform_sig_rx =-719;
5603: waveform_sig_rx =-545;
5604: waveform_sig_rx =-1015;
5605: waveform_sig_rx =-559;
5606: waveform_sig_rx =-691;
5607: waveform_sig_rx =-955;
5608: waveform_sig_rx =-575;
5609: waveform_sig_rx =-716;
5610: waveform_sig_rx =-931;
5611: waveform_sig_rx =-684;
5612: waveform_sig_rx =-688;
5613: waveform_sig_rx =-923;
5614: waveform_sig_rx =-780;
5615: waveform_sig_rx =-653;
5616: waveform_sig_rx =-884;
5617: waveform_sig_rx =-928;
5618: waveform_sig_rx =-590;
5619: waveform_sig_rx =-867;
5620: waveform_sig_rx =-944;
5621: waveform_sig_rx =-740;
5622: waveform_sig_rx =-732;
5623: waveform_sig_rx =-1034;
5624: waveform_sig_rx =-738;
5625: waveform_sig_rx =-748;
5626: waveform_sig_rx =-978;
5627: waveform_sig_rx =-870;
5628: waveform_sig_rx =-737;
5629: waveform_sig_rx =-879;
5630: waveform_sig_rx =-1011;
5631: waveform_sig_rx =-749;
5632: waveform_sig_rx =-824;
5633: waveform_sig_rx =-1081;
5634: waveform_sig_rx =-786;
5635: waveform_sig_rx =-760;
5636: waveform_sig_rx =-1111;
5637: waveform_sig_rx =-769;
5638: waveform_sig_rx =-996;
5639: waveform_sig_rx =-887;
5640: waveform_sig_rx =-898;
5641: waveform_sig_rx =-874;
5642: waveform_sig_rx =-1018;
5643: waveform_sig_rx =-897;
5644: waveform_sig_rx =-827;
5645: waveform_sig_rx =-1166;
5646: waveform_sig_rx =-784;
5647: waveform_sig_rx =-930;
5648: waveform_sig_rx =-1110;
5649: waveform_sig_rx =-827;
5650: waveform_sig_rx =-878;
5651: waveform_sig_rx =-1137;
5652: waveform_sig_rx =-898;
5653: waveform_sig_rx =-834;
5654: waveform_sig_rx =-1158;
5655: waveform_sig_rx =-965;
5656: waveform_sig_rx =-849;
5657: waveform_sig_rx =-1129;
5658: waveform_sig_rx =-1099;
5659: waveform_sig_rx =-795;
5660: waveform_sig_rx =-1091;
5661: waveform_sig_rx =-1091;
5662: waveform_sig_rx =-931;
5663: waveform_sig_rx =-948;
5664: waveform_sig_rx =-1185;
5665: waveform_sig_rx =-940;
5666: waveform_sig_rx =-960;
5667: waveform_sig_rx =-1143;
5668: waveform_sig_rx =-1086;
5669: waveform_sig_rx =-896;
5670: waveform_sig_rx =-1055;
5671: waveform_sig_rx =-1220;
5672: waveform_sig_rx =-843;
5673: waveform_sig_rx =-1051;
5674: waveform_sig_rx =-1253;
5675: waveform_sig_rx =-904;
5676: waveform_sig_rx =-1012;
5677: waveform_sig_rx =-1238;
5678: waveform_sig_rx =-924;
5679: waveform_sig_rx =-1212;
5680: waveform_sig_rx =-985;
5681: waveform_sig_rx =-1115;
5682: waveform_sig_rx =-1053;
5683: waveform_sig_rx =-1148;
5684: waveform_sig_rx =-1091;
5685: waveform_sig_rx =-982;
5686: waveform_sig_rx =-1273;
5687: waveform_sig_rx =-970;
5688: waveform_sig_rx =-1053;
5689: waveform_sig_rx =-1286;
5690: waveform_sig_rx =-988;
5691: waveform_sig_rx =-1008;
5692: waveform_sig_rx =-1342;
5693: waveform_sig_rx =-1001;
5694: waveform_sig_rx =-983;
5695: waveform_sig_rx =-1342;
5696: waveform_sig_rx =-1042;
5697: waveform_sig_rx =-980;
5698: waveform_sig_rx =-1268;
5699: waveform_sig_rx =-1156;
5700: waveform_sig_rx =-934;
5701: waveform_sig_rx =-1216;
5702: waveform_sig_rx =-1170;
5703: waveform_sig_rx =-1062;
5704: waveform_sig_rx =-1051;
5705: waveform_sig_rx =-1265;
5706: waveform_sig_rx =-1082;
5707: waveform_sig_rx =-1005;
5708: waveform_sig_rx =-1246;
5709: waveform_sig_rx =-1212;
5710: waveform_sig_rx =-930;
5711: waveform_sig_rx =-1242;
5712: waveform_sig_rx =-1280;
5713: waveform_sig_rx =-933;
5714: waveform_sig_rx =-1242;
5715: waveform_sig_rx =-1260;
5716: waveform_sig_rx =-1032;
5717: waveform_sig_rx =-1112;
5718: waveform_sig_rx =-1252;
5719: waveform_sig_rx =-1076;
5720: waveform_sig_rx =-1237;
5721: waveform_sig_rx =-1056;
5722: waveform_sig_rx =-1217;
5723: waveform_sig_rx =-1062;
5724: waveform_sig_rx =-1256;
5725: waveform_sig_rx =-1142;
5726: waveform_sig_rx =-1043;
5727: waveform_sig_rx =-1366;
5728: waveform_sig_rx =-1028;
5729: waveform_sig_rx =-1090;
5730: waveform_sig_rx =-1367;
5731: waveform_sig_rx =-1029;
5732: waveform_sig_rx =-1035;
5733: waveform_sig_rx =-1445;
5734: waveform_sig_rx =-991;
5735: waveform_sig_rx =-1070;
5736: waveform_sig_rx =-1420;
5737: waveform_sig_rx =-1010;
5738: waveform_sig_rx =-1116;
5739: waveform_sig_rx =-1299;
5740: waveform_sig_rx =-1170;
5741: waveform_sig_rx =-1061;
5742: waveform_sig_rx =-1205;
5743: waveform_sig_rx =-1241;
5744: waveform_sig_rx =-1104;
5745: waveform_sig_rx =-1045;
5746: waveform_sig_rx =-1365;
5747: waveform_sig_rx =-1070;
5748: waveform_sig_rx =-1044;
5749: waveform_sig_rx =-1321;
5750: waveform_sig_rx =-1172;
5751: waveform_sig_rx =-970;
5752: waveform_sig_rx =-1281;
5753: waveform_sig_rx =-1236;
5754: waveform_sig_rx =-983;
5755: waveform_sig_rx =-1232;
5756: waveform_sig_rx =-1226;
5757: waveform_sig_rx =-1058;
5758: waveform_sig_rx =-1099;
5759: waveform_sig_rx =-1260;
5760: waveform_sig_rx =-1118;
5761: waveform_sig_rx =-1196;
5762: waveform_sig_rx =-1069;
5763: waveform_sig_rx =-1246;
5764: waveform_sig_rx =-1020;
5765: waveform_sig_rx =-1280;
5766: waveform_sig_rx =-1104;
5767: waveform_sig_rx =-1025;
5768: waveform_sig_rx =-1380;
5769: waveform_sig_rx =-970;
5770: waveform_sig_rx =-1109;
5771: waveform_sig_rx =-1354;
5772: waveform_sig_rx =-940;
5773: waveform_sig_rx =-1084;
5774: waveform_sig_rx =-1383;
5775: waveform_sig_rx =-914;
5776: waveform_sig_rx =-1103;
5777: waveform_sig_rx =-1325;
5778: waveform_sig_rx =-964;
5779: waveform_sig_rx =-1104;
5780: waveform_sig_rx =-1191;
5781: waveform_sig_rx =-1148;
5782: waveform_sig_rx =-1003;
5783: waveform_sig_rx =-1124;
5784: waveform_sig_rx =-1239;
5785: waveform_sig_rx =-993;
5786: waveform_sig_rx =-999;
5787: waveform_sig_rx =-1330;
5788: waveform_sig_rx =-941;
5789: waveform_sig_rx =-1032;
5790: waveform_sig_rx =-1236;
5791: waveform_sig_rx =-1041;
5792: waveform_sig_rx =-938;
5793: waveform_sig_rx =-1195;
5794: waveform_sig_rx =-1134;
5795: waveform_sig_rx =-917;
5796: waveform_sig_rx =-1119;
5797: waveform_sig_rx =-1159;
5798: waveform_sig_rx =-980;
5799: waveform_sig_rx =-964;
5800: waveform_sig_rx =-1201;
5801: waveform_sig_rx =-996;
5802: waveform_sig_rx =-1085;
5803: waveform_sig_rx =-1005;
5804: waveform_sig_rx =-1089;
5805: waveform_sig_rx =-918;
5806: waveform_sig_rx =-1230;
5807: waveform_sig_rx =-915;
5808: waveform_sig_rx =-970;
5809: waveform_sig_rx =-1269;
5810: waveform_sig_rx =-801;
5811: waveform_sig_rx =-1069;
5812: waveform_sig_rx =-1183;
5813: waveform_sig_rx =-803;
5814: waveform_sig_rx =-1038;
5815: waveform_sig_rx =-1220;
5816: waveform_sig_rx =-801;
5817: waveform_sig_rx =-1011;
5818: waveform_sig_rx =-1131;
5819: waveform_sig_rx =-891;
5820: waveform_sig_rx =-938;
5821: waveform_sig_rx =-1077;
5822: waveform_sig_rx =-1057;
5823: waveform_sig_rx =-811;
5824: waveform_sig_rx =-1041;
5825: waveform_sig_rx =-1114;
5826: waveform_sig_rx =-821;
5827: waveform_sig_rx =-927;
5828: waveform_sig_rx =-1173;
5829: waveform_sig_rx =-787;
5830: waveform_sig_rx =-942;
5831: waveform_sig_rx =-1081;
5832: waveform_sig_rx =-918;
5833: waveform_sig_rx =-836;
5834: waveform_sig_rx =-1009;
5835: waveform_sig_rx =-1013;
5836: waveform_sig_rx =-767;
5837: waveform_sig_rx =-941;
5838: waveform_sig_rx =-1071;
5839: waveform_sig_rx =-763;
5840: waveform_sig_rx =-855;
5841: waveform_sig_rx =-1080;
5842: waveform_sig_rx =-767;
5843: waveform_sig_rx =-992;
5844: waveform_sig_rx =-846;
5845: waveform_sig_rx =-919;
5846: waveform_sig_rx =-810;
5847: waveform_sig_rx =-1038;
5848: waveform_sig_rx =-743;
5849: waveform_sig_rx =-855;
5850: waveform_sig_rx =-1065;
5851: waveform_sig_rx =-645;
5852: waveform_sig_rx =-922;
5853: waveform_sig_rx =-985;
5854: waveform_sig_rx =-637;
5855: waveform_sig_rx =-886;
5856: waveform_sig_rx =-1003;
5857: waveform_sig_rx =-683;
5858: waveform_sig_rx =-814;
5859: waveform_sig_rx =-952;
5860: waveform_sig_rx =-750;
5861: waveform_sig_rx =-687;
5862: waveform_sig_rx =-972;
5863: waveform_sig_rx =-842;
5864: waveform_sig_rx =-579;
5865: waveform_sig_rx =-944;
5866: waveform_sig_rx =-834;
5867: waveform_sig_rx =-629;
5868: waveform_sig_rx =-782;
5869: waveform_sig_rx =-894;
5870: waveform_sig_rx =-652;
5871: waveform_sig_rx =-704;
5872: waveform_sig_rx =-852;
5873: waveform_sig_rx =-733;
5874: waveform_sig_rx =-585;
5875: waveform_sig_rx =-846;
5876: waveform_sig_rx =-817;
5877: waveform_sig_rx =-530;
5878: waveform_sig_rx =-771;
5879: waveform_sig_rx =-852;
5880: waveform_sig_rx =-534;
5881: waveform_sig_rx =-684;
5882: waveform_sig_rx =-840;
5883: waveform_sig_rx =-553;
5884: waveform_sig_rx =-809;
5885: waveform_sig_rx =-585;
5886: waveform_sig_rx =-696;
5887: waveform_sig_rx =-615;
5888: waveform_sig_rx =-783;
5889: waveform_sig_rx =-512;
5890: waveform_sig_rx =-658;
5891: waveform_sig_rx =-774;
5892: waveform_sig_rx =-452;
5893: waveform_sig_rx =-679;
5894: waveform_sig_rx =-720;
5895: waveform_sig_rx =-463;
5896: waveform_sig_rx =-587;
5897: waveform_sig_rx =-798;
5898: waveform_sig_rx =-427;
5899: waveform_sig_rx =-540;
5900: waveform_sig_rx =-780;
5901: waveform_sig_rx =-449;
5902: waveform_sig_rx =-467;
5903: waveform_sig_rx =-754;
5904: waveform_sig_rx =-522;
5905: waveform_sig_rx =-407;
5906: waveform_sig_rx =-665;
5907: waveform_sig_rx =-561;
5908: waveform_sig_rx =-442;
5909: waveform_sig_rx =-500;
5910: waveform_sig_rx =-658;
5911: waveform_sig_rx =-400;
5912: waveform_sig_rx =-444;
5913: waveform_sig_rx =-629;
5914: waveform_sig_rx =-478;
5915: waveform_sig_rx =-330;
5916: waveform_sig_rx =-609;
5917: waveform_sig_rx =-541;
5918: waveform_sig_rx =-279;
5919: waveform_sig_rx =-570;
5920: waveform_sig_rx =-578;
5921: waveform_sig_rx =-247;
5922: waveform_sig_rx =-486;
5923: waveform_sig_rx =-514;
5924: waveform_sig_rx =-311;
5925: waveform_sig_rx =-586;
5926: waveform_sig_rx =-274;
5927: waveform_sig_rx =-518;
5928: waveform_sig_rx =-319;
5929: waveform_sig_rx =-492;
5930: waveform_sig_rx =-317;
5931: waveform_sig_rx =-326;
5932: waveform_sig_rx =-536;
5933: waveform_sig_rx =-209;
5934: waveform_sig_rx =-364;
5935: waveform_sig_rx =-546;
5936: waveform_sig_rx =-128;
5937: waveform_sig_rx =-346;
5938: waveform_sig_rx =-573;
5939: waveform_sig_rx =-74;
5940: waveform_sig_rx =-361;
5941: waveform_sig_rx =-479;
5942: waveform_sig_rx =-161;
5943: waveform_sig_rx =-270;
5944: waveform_sig_rx =-458;
5945: waveform_sig_rx =-241;
5946: waveform_sig_rx =-170;
5947: waveform_sig_rx =-373;
5948: waveform_sig_rx =-305;
5949: waveform_sig_rx =-156;
5950: waveform_sig_rx =-218;
5951: waveform_sig_rx =-383;
5952: waveform_sig_rx =-107;
5953: waveform_sig_rx =-157;
5954: waveform_sig_rx =-374;
5955: waveform_sig_rx =-176;
5956: waveform_sig_rx =-21;
5957: waveform_sig_rx =-382;
5958: waveform_sig_rx =-200;
5959: waveform_sig_rx =6;
5960: waveform_sig_rx =-320;
5961: waveform_sig_rx =-198;
5962: waveform_sig_rx =-30;
5963: waveform_sig_rx =-200;
5964: waveform_sig_rx =-173;
5965: waveform_sig_rx =-121;
5966: waveform_sig_rx =-192;
5967: waveform_sig_rx =-8;
5968: waveform_sig_rx =-242;
5969: waveform_sig_rx =69;
5970: waveform_sig_rx =-292;
5971: waveform_sig_rx =40;
5972: waveform_sig_rx =-42;
5973: waveform_sig_rx =-317;
5974: waveform_sig_rx =178;
5975: waveform_sig_rx =-162;
5976: waveform_sig_rx =-247;
5977: waveform_sig_rx =220;
5978: waveform_sig_rx =-140;
5979: waveform_sig_rx =-196;
5980: waveform_sig_rx =199;
5981: waveform_sig_rx =-78;
5982: waveform_sig_rx =-175;
5983: waveform_sig_rx =104;
5984: waveform_sig_rx =24;
5985: waveform_sig_rx =-188;
5986: waveform_sig_rx =82;
5987: waveform_sig_rx =85;
5988: waveform_sig_rx =-67;
5989: waveform_sig_rx =-23;
5990: waveform_sig_rx =116;
5991: waveform_sig_rx =126;
5992: waveform_sig_rx =-179;
5993: waveform_sig_rx =237;
5994: waveform_sig_rx =139;
5995: waveform_sig_rx =-154;
5996: waveform_sig_rx =244;
5997: waveform_sig_rx =156;
5998: waveform_sig_rx =-42;
5999: waveform_sig_rx =157;
6000: waveform_sig_rx =208;
6001: waveform_sig_rx =99;
6002: waveform_sig_rx =30;
6003: waveform_sig_rx =283;
6004: waveform_sig_rx =177;
6005: waveform_sig_rx =30;
6006: waveform_sig_rx =242;
6007: waveform_sig_rx =101;
6008: waveform_sig_rx =235;
6009: waveform_sig_rx =134;
6010: waveform_sig_rx =308;
6011: waveform_sig_rx =-36;
6012: waveform_sig_rx =381;
6013: waveform_sig_rx =178;
6014: waveform_sig_rx =4;
6015: waveform_sig_rx =494;
6016: waveform_sig_rx =88;
6017: waveform_sig_rx =102;
6018: waveform_sig_rx =533;
6019: waveform_sig_rx =114;
6020: waveform_sig_rx =150;
6021: waveform_sig_rx =496;
6022: waveform_sig_rx =185;
6023: waveform_sig_rx =213;
6024: waveform_sig_rx =382;
6025: waveform_sig_rx =329;
6026: waveform_sig_rx =159;
6027: waveform_sig_rx =326;
6028: waveform_sig_rx =414;
6029: waveform_sig_rx =224;
6030: waveform_sig_rx =208;
6031: waveform_sig_rx =488;
6032: waveform_sig_rx =337;
6033: waveform_sig_rx =146;
6034: waveform_sig_rx =605;
6035: waveform_sig_rx =313;
6036: waveform_sig_rx =216;
6037: waveform_sig_rx =497;
6038: waveform_sig_rx =412;
6039: waveform_sig_rx =314;
6040: waveform_sig_rx =347;
6041: waveform_sig_rx =533;
6042: waveform_sig_rx =371;
6043: waveform_sig_rx =255;
6044: waveform_sig_rx =628;
6045: waveform_sig_rx =381;
6046: waveform_sig_rx =309;
6047: waveform_sig_rx =556;
6048: waveform_sig_rx =337;
6049: waveform_sig_rx =542;
6050: waveform_sig_rx =411;
6051: waveform_sig_rx =542;
6052: waveform_sig_rx =281;
6053: waveform_sig_rx =665;
6054: waveform_sig_rx =407;
6055: waveform_sig_rx =337;
6056: waveform_sig_rx =755;
6057: waveform_sig_rx =323;
6058: waveform_sig_rx =440;
6059: waveform_sig_rx =754;
6060: waveform_sig_rx =349;
6061: waveform_sig_rx =453;
6062: waveform_sig_rx =713;
6063: waveform_sig_rx =465;
6064: waveform_sig_rx =483;
6065: waveform_sig_rx =600;
6066: waveform_sig_rx =673;
6067: waveform_sig_rx =366;
6068: waveform_sig_rx =593;
6069: waveform_sig_rx =762;
6070: waveform_sig_rx =408;
6071: waveform_sig_rx =561;
6072: waveform_sig_rx =750;
6073: waveform_sig_rx =524;
6074: waveform_sig_rx =510;
6075: waveform_sig_rx =791;
6076: waveform_sig_rx =580;
6077: waveform_sig_rx =532;
6078: waveform_sig_rx =699;
6079: waveform_sig_rx =742;
6080: waveform_sig_rx =531;
6081: waveform_sig_rx =609;
6082: waveform_sig_rx =841;
6083: waveform_sig_rx =578;
6084: waveform_sig_rx =546;
6085: waveform_sig_rx =908;
6086: waveform_sig_rx =590;
6087: waveform_sig_rx =599;
6088: waveform_sig_rx =816;
6089: waveform_sig_rx =571;
6090: waveform_sig_rx =799;
6091: waveform_sig_rx =673;
6092: waveform_sig_rx =749;
6093: waveform_sig_rx =576;
6094: waveform_sig_rx =919;
6095: waveform_sig_rx =619;
6096: waveform_sig_rx =666;
6097: waveform_sig_rx =928;
6098: waveform_sig_rx =595;
6099: waveform_sig_rx =724;
6100: waveform_sig_rx =925;
6101: waveform_sig_rx =679;
6102: waveform_sig_rx =666;
6103: waveform_sig_rx =946;
6104: waveform_sig_rx =746;
6105: waveform_sig_rx =649;
6106: waveform_sig_rx =913;
6107: waveform_sig_rx =889;
6108: waveform_sig_rx =578;
6109: waveform_sig_rx =915;
6110: waveform_sig_rx =921;
6111: waveform_sig_rx =655;
6112: waveform_sig_rx =836;
6113: waveform_sig_rx =948;
6114: waveform_sig_rx =759;
6115: waveform_sig_rx =757;
6116: waveform_sig_rx =961;
6117: waveform_sig_rx =832;
6118: waveform_sig_rx =748;
6119: waveform_sig_rx =895;
6120: waveform_sig_rx =999;
6121: waveform_sig_rx =696;
6122: waveform_sig_rx =829;
6123: waveform_sig_rx =1083;
6124: waveform_sig_rx =705;
6125: waveform_sig_rx =834;
6126: waveform_sig_rx =1106;
6127: waveform_sig_rx =759;
6128: waveform_sig_rx =890;
6129: waveform_sig_rx =963;
6130: waveform_sig_rx =802;
6131: waveform_sig_rx =1053;
6132: waveform_sig_rx =850;
6133: waveform_sig_rx =985;
6134: waveform_sig_rx =787;
6135: waveform_sig_rx =1079;
6136: waveform_sig_rx =843;
6137: waveform_sig_rx =865;
6138: waveform_sig_rx =1104;
6139: waveform_sig_rx =833;
6140: waveform_sig_rx =877;
6141: waveform_sig_rx =1156;
6142: waveform_sig_rx =892;
6143: waveform_sig_rx =799;
6144: waveform_sig_rx =1207;
6145: waveform_sig_rx =898;
6146: waveform_sig_rx =815;
6147: waveform_sig_rx =1164;
6148: waveform_sig_rx =1005;
6149: waveform_sig_rx =780;
6150: waveform_sig_rx =1123;
6151: waveform_sig_rx =1019;
6152: waveform_sig_rx =872;
6153: waveform_sig_rx =998;
6154: waveform_sig_rx =1100;
6155: waveform_sig_rx =976;
6156: waveform_sig_rx =897;
6157: waveform_sig_rx =1148;
6158: waveform_sig_rx =1038;
6159: waveform_sig_rx =867;
6160: waveform_sig_rx =1104;
6161: waveform_sig_rx =1165;
6162: waveform_sig_rx =825;
6163: waveform_sig_rx =1092;
6164: waveform_sig_rx =1214;
6165: waveform_sig_rx =853;
6166: waveform_sig_rx =1047;
6167: waveform_sig_rx =1219;
6168: waveform_sig_rx =918;
6169: waveform_sig_rx =1061;
6170: waveform_sig_rx =1059;
6171: waveform_sig_rx =994;
6172: waveform_sig_rx =1174;
6173: waveform_sig_rx =991;
6174: waveform_sig_rx =1175;
6175: waveform_sig_rx =897;
6176: waveform_sig_rx =1237;
6177: waveform_sig_rx =1001;
6178: waveform_sig_rx =974;
6179: waveform_sig_rx =1274;
6180: waveform_sig_rx =971;
6181: waveform_sig_rx =981;
6182: waveform_sig_rx =1350;
6183: waveform_sig_rx =962;
6184: waveform_sig_rx =929;
6185: waveform_sig_rx =1369;
6186: waveform_sig_rx =931;
6187: waveform_sig_rx =1008;
6188: waveform_sig_rx =1286;
6189: waveform_sig_rx =1055;
6190: waveform_sig_rx =984;
6191: waveform_sig_rx =1226;
6192: waveform_sig_rx =1148;
6193: waveform_sig_rx =1042;
6194: waveform_sig_rx =1067;
6195: waveform_sig_rx =1254;
6196: waveform_sig_rx =1081;
6197: waveform_sig_rx =981;
6198: waveform_sig_rx =1325;
6199: waveform_sig_rx =1089;
6200: waveform_sig_rx =956;
6201: waveform_sig_rx =1267;
6202: waveform_sig_rx =1198;
6203: waveform_sig_rx =918;
6204: waveform_sig_rx =1199;
6205: waveform_sig_rx =1249;
6206: waveform_sig_rx =989;
6207: waveform_sig_rx =1149;
6208: waveform_sig_rx =1276;
6209: waveform_sig_rx =1076;
6210: waveform_sig_rx =1140;
6211: waveform_sig_rx =1147;
6212: waveform_sig_rx =1142;
6213: waveform_sig_rx =1191;
6214: waveform_sig_rx =1087;
6215: waveform_sig_rx =1257;
6216: waveform_sig_rx =939;
6217: waveform_sig_rx =1365;
6218: waveform_sig_rx =1036;
6219: waveform_sig_rx =1035;
6220: waveform_sig_rx =1396;
6221: waveform_sig_rx =960;
6222: waveform_sig_rx =1089;
6223: waveform_sig_rx =1414;
6224: waveform_sig_rx =949;
6225: waveform_sig_rx =1091;
6226: waveform_sig_rx =1414;
6227: waveform_sig_rx =962;
6228: waveform_sig_rx =1140;
6229: waveform_sig_rx =1284;
6230: waveform_sig_rx =1128;
6231: waveform_sig_rx =1034;
6232: waveform_sig_rx =1234;
6233: waveform_sig_rx =1247;
6234: waveform_sig_rx =1053;
6235: waveform_sig_rx =1103;
6236: waveform_sig_rx =1331;
6237: waveform_sig_rx =1047;
6238: waveform_sig_rx =1037;
6239: waveform_sig_rx =1345;
6240: waveform_sig_rx =1088;
6241: waveform_sig_rx =1018;
6242: waveform_sig_rx =1302;
6243: waveform_sig_rx =1184;
6244: waveform_sig_rx =976;
6245: waveform_sig_rx =1253;
6246: waveform_sig_rx =1217;
6247: waveform_sig_rx =1049;
6248: waveform_sig_rx =1119;
6249: waveform_sig_rx =1280;
6250: waveform_sig_rx =1105;
6251: waveform_sig_rx =1077;
6252: waveform_sig_rx =1194;
6253: waveform_sig_rx =1119;
6254: waveform_sig_rx =1153;
6255: waveform_sig_rx =1169;
6256: waveform_sig_rx =1171;
6257: waveform_sig_rx =974;
6258: waveform_sig_rx =1409;
6259: waveform_sig_rx =954;
6260: waveform_sig_rx =1123;
6261: waveform_sig_rx =1360;
6262: waveform_sig_rx =930;
6263: waveform_sig_rx =1141;
6264: waveform_sig_rx =1338;
6265: waveform_sig_rx =946;
6266: waveform_sig_rx =1081;
6267: waveform_sig_rx =1343;
6268: waveform_sig_rx =952;
6269: waveform_sig_rx =1126;
6270: waveform_sig_rx =1228;
6271: waveform_sig_rx =1128;
6272: waveform_sig_rx =988;
6273: waveform_sig_rx =1183;
6274: waveform_sig_rx =1212;
6275: waveform_sig_rx =975;
6276: waveform_sig_rx =1098;
6277: waveform_sig_rx =1320;
6278: waveform_sig_rx =958;
6279: waveform_sig_rx =1090;
6280: waveform_sig_rx =1294;
6281: waveform_sig_rx =1008;
6282: waveform_sig_rx =1047;
6283: waveform_sig_rx =1182;
6284: waveform_sig_rx =1153;
6285: waveform_sig_rx =969;
6286: waveform_sig_rx =1164;
6287: waveform_sig_rx =1239;
6288: waveform_sig_rx =958;
6289: waveform_sig_rx =1047;
6290: waveform_sig_rx =1285;
6291: waveform_sig_rx =964;
6292: waveform_sig_rx =1075;
6293: waveform_sig_rx =1137;
6294: waveform_sig_rx =1007;
6295: waveform_sig_rx =1115;
6296: waveform_sig_rx =1089;
6297: waveform_sig_rx =1062;
6298: waveform_sig_rx =956;
6299: waveform_sig_rx =1288;
6300: waveform_sig_rx =852;
6301: waveform_sig_rx =1094;
6302: waveform_sig_rx =1203;
6303: waveform_sig_rx =866;
6304: waveform_sig_rx =1078;
6305: waveform_sig_rx =1215;
6306: waveform_sig_rx =900;
6307: waveform_sig_rx =1012;
6308: waveform_sig_rx =1226;
6309: waveform_sig_rx =891;
6310: waveform_sig_rx =1011;
6311: waveform_sig_rx =1127;
6312: waveform_sig_rx =1040;
6313: waveform_sig_rx =824;
6314: waveform_sig_rx =1154;
6315: waveform_sig_rx =1102;
6316: waveform_sig_rx =832;
6317: waveform_sig_rx =1055;
6318: waveform_sig_rx =1158;
6319: waveform_sig_rx =831;
6320: waveform_sig_rx =1020;
6321: waveform_sig_rx =1103;
6322: waveform_sig_rx =946;
6323: waveform_sig_rx =904;
6324: waveform_sig_rx =1034;
6325: waveform_sig_rx =1073;
6326: waveform_sig_rx =766;
6327: waveform_sig_rx =1058;
6328: waveform_sig_rx =1092;
6329: waveform_sig_rx =790;
6330: waveform_sig_rx =985;
6331: waveform_sig_rx =1132;
6332: waveform_sig_rx =818;
6333: waveform_sig_rx =983;
6334: waveform_sig_rx =962;
6335: waveform_sig_rx =885;
6336: waveform_sig_rx =995;
6337: waveform_sig_rx =913;
6338: waveform_sig_rx =919;
6339: waveform_sig_rx =837;
6340: waveform_sig_rx =1100;
6341: waveform_sig_rx =728;
6342: waveform_sig_rx =936;
6343: waveform_sig_rx =1016;
6344: waveform_sig_rx =757;
6345: waveform_sig_rx =905;
6346: waveform_sig_rx =1054;
6347: waveform_sig_rx =760;
6348: waveform_sig_rx =807;
6349: waveform_sig_rx =1112;
6350: waveform_sig_rx =724;
6351: waveform_sig_rx =796;
6352: waveform_sig_rx =1050;
6353: waveform_sig_rx =808;
6354: waveform_sig_rx =686;
6355: waveform_sig_rx =1034;
6356: waveform_sig_rx =831;
6357: waveform_sig_rx =731;
6358: waveform_sig_rx =867;
6359: waveform_sig_rx =927;
6360: waveform_sig_rx =718;
6361: waveform_sig_rx =782;
6362: waveform_sig_rx =949;
6363: waveform_sig_rx =756;
6364: waveform_sig_rx =677;
6365: waveform_sig_rx =927;
6366: waveform_sig_rx =846;
6367: waveform_sig_rx =586;
6368: waveform_sig_rx =886;
6369: waveform_sig_rx =900;
6370: waveform_sig_rx =563;
6371: waveform_sig_rx =811;
6372: waveform_sig_rx =929;
6373: waveform_sig_rx =571;
6374: waveform_sig_rx =840;
6375: waveform_sig_rx =687;
6376: waveform_sig_rx =708;
6377: waveform_sig_rx =812;
6378: waveform_sig_rx =661;
6379: waveform_sig_rx =778;
6380: waveform_sig_rx =596;
6381: waveform_sig_rx =874;
6382: waveform_sig_rx =584;
6383: waveform_sig_rx =671;
6384: waveform_sig_rx =851;
6385: waveform_sig_rx =502;
6386: waveform_sig_rx =644;
6387: waveform_sig_rx =876;
6388: waveform_sig_rx =449;
6389: waveform_sig_rx =625;
6390: waveform_sig_rx =866;
6391: waveform_sig_rx =437;
6392: waveform_sig_rx =637;
6393: waveform_sig_rx =783;
6394: waveform_sig_rx =569;
6395: waveform_sig_rx =483;
6396: waveform_sig_rx =787;
6397: waveform_sig_rx =584;
6398: waveform_sig_rx =516;
6399: waveform_sig_rx =620;
6400: waveform_sig_rx =703;
6401: waveform_sig_rx =500;
6402: waveform_sig_rx =518;
6403: waveform_sig_rx =738;
6404: waveform_sig_rx =514;
6405: waveform_sig_rx =413;
6406: waveform_sig_rx =743;
6407: waveform_sig_rx =589;
6408: waveform_sig_rx =335;
6409: waveform_sig_rx =708;
6410: waveform_sig_rx =580;
6411: waveform_sig_rx =345;
6412: waveform_sig_rx =596;
6413: waveform_sig_rx =608;
6414: waveform_sig_rx =382;
6415: waveform_sig_rx =582;
6416: waveform_sig_rx =419;
6417: waveform_sig_rx =530;
6418: waveform_sig_rx =470;
6419: waveform_sig_rx =443;
6420: waveform_sig_rx =521;
6421: waveform_sig_rx =279;
6422: waveform_sig_rx =683;
6423: waveform_sig_rx =259;
6424: waveform_sig_rx =412;
6425: waveform_sig_rx =645;
6426: waveform_sig_rx =162;
6427: waveform_sig_rx =479;
6428: waveform_sig_rx =597;
6429: waveform_sig_rx =151;
6430: waveform_sig_rx =420;
6431: waveform_sig_rx =554;
6432: waveform_sig_rx =189;
6433: waveform_sig_rx =358;
6434: waveform_sig_rx =507;
6435: waveform_sig_rx =284;
6436: waveform_sig_rx =223;
6437: waveform_sig_rx =528;
6438: waveform_sig_rx =280;
6439: waveform_sig_rx =281;
6440: waveform_sig_rx =298;
6441: waveform_sig_rx =448;
6442: waveform_sig_rx =199;
6443: waveform_sig_rx =206;
6444: waveform_sig_rx =534;
6445: waveform_sig_rx =156;
6446: waveform_sig_rx =165;
6447: waveform_sig_rx =512;
6448: waveform_sig_rx =172;
6449: waveform_sig_rx =155;
6450: waveform_sig_rx =362;
6451: waveform_sig_rx =253;
6452: waveform_sig_rx =142;
6453: waveform_sig_rx =201;
6454: waveform_sig_rx =378;
6455: waveform_sig_rx =71;
6456: waveform_sig_rx =221;
6457: waveform_sig_rx =196;
6458: waveform_sig_rx =200;
6459: waveform_sig_rx =165;
6460: waveform_sig_rx =223;
6461: waveform_sig_rx =146;
6462: waveform_sig_rx =30;
6463: waveform_sig_rx =393;
6464: waveform_sig_rx =-95;
6465: waveform_sig_rx =183;
6466: waveform_sig_rx =301;
6467: waveform_sig_rx =-137;
6468: waveform_sig_rx =202;
6469: waveform_sig_rx =267;
6470: waveform_sig_rx =-146;
6471: waveform_sig_rx =158;
6472: waveform_sig_rx =232;
6473: waveform_sig_rx =-137;
6474: waveform_sig_rx =118;
6475: waveform_sig_rx =149;
6476: waveform_sig_rx =4;
6477: waveform_sig_rx =-79;
6478: waveform_sig_rx =140;
6479: waveform_sig_rx =49;
6480: waveform_sig_rx =-97;
6481: waveform_sig_rx =5;
6482: waveform_sig_rx =215;
6483: waveform_sig_rx =-220;
6484: waveform_sig_rx =-1;
6485: waveform_sig_rx =183;
6486: waveform_sig_rx =-203;
6487: waveform_sig_rx =-39;
6488: waveform_sig_rx =77;
6489: waveform_sig_rx =-73;
6490: waveform_sig_rx =-139;
6491: waveform_sig_rx =-21;
6492: waveform_sig_rx =17;
6493: waveform_sig_rx =-236;
6494: waveform_sig_rx =-63;
6495: waveform_sig_rx =98;
6496: waveform_sig_rx =-281;
6497: waveform_sig_rx =-22;
6498: waveform_sig_rx =-134;
6499: waveform_sig_rx =-106;
6500: waveform_sig_rx =-110;
6501: waveform_sig_rx =-96;
6502: waveform_sig_rx =-168;
6503: waveform_sig_rx =-242;
6504: waveform_sig_rx =69;
6505: waveform_sig_rx =-424;
6506: waveform_sig_rx =-80;
6507: waveform_sig_rx =-43;
6508: waveform_sig_rx =-466;
6509: waveform_sig_rx =-37;
6510: waveform_sig_rx =-112;
6511: waveform_sig_rx =-428;
6512: waveform_sig_rx =-115;
6513: waveform_sig_rx =-136;
6514: waveform_sig_rx =-347;
6515: waveform_sig_rx =-239;
6516: waveform_sig_rx =-138;
6517: waveform_sig_rx =-259;
6518: waveform_sig_rx =-452;
6519: waveform_sig_rx =-58;
6520: waveform_sig_rx =-302;
6521: waveform_sig_rx =-443;
6522: waveform_sig_rx =-204;
6523: waveform_sig_rx =-179;
6524: waveform_sig_rx =-466;
6525: waveform_sig_rx =-280;
6526: waveform_sig_rx =-200;
6527: waveform_sig_rx =-449;
6528: waveform_sig_rx =-379;
6529: waveform_sig_rx =-222;
6530: waveform_sig_rx =-357;
6531: waveform_sig_rx =-521;
6532: waveform_sig_rx =-277;
6533: waveform_sig_rx =-274;
6534: waveform_sig_rx =-572;
6535: waveform_sig_rx =-339;
6536: waveform_sig_rx =-224;
6537: waveform_sig_rx =-602;
6538: waveform_sig_rx =-302;
6539: waveform_sig_rx =-477;
6540: waveform_sig_rx =-412;
6541: waveform_sig_rx =-392;
6542: waveform_sig_rx =-395;
6543: waveform_sig_rx =-514;
6544: waveform_sig_rx =-485;
6545: waveform_sig_rx =-285;
6546: waveform_sig_rx =-703;
6547: waveform_sig_rx =-336;
6548: waveform_sig_rx =-426;
6549: waveform_sig_rx =-672;
6550: waveform_sig_rx =-365;
6551: waveform_sig_rx =-436;
6552: waveform_sig_rx =-653;
6553: waveform_sig_rx =-478;
6554: waveform_sig_rx =-376;
6555: waveform_sig_rx =-656;
6556: waveform_sig_rx =-578;
6557: waveform_sig_rx =-340;
6558: waveform_sig_rx =-613;
6559: waveform_sig_rx =-716;
6560: waveform_sig_rx =-289;
6561: waveform_sig_rx =-654;
6562: waveform_sig_rx =-638;
6563: waveform_sig_rx =-498;
6564: waveform_sig_rx =-494;
6565: waveform_sig_rx =-705;
6566: waveform_sig_rx =-578;
6567: waveform_sig_rx =-469;
6568: waveform_sig_rx =-696;
6569: waveform_sig_rx =-667;
6570: waveform_sig_rx =-458;
6571: waveform_sig_rx =-622;
6572: waveform_sig_rx =-798;
6573: waveform_sig_rx =-513;
6574: waveform_sig_rx =-565;
6575: waveform_sig_rx =-857;
6576: waveform_sig_rx =-543;
6577: waveform_sig_rx =-528;
6578: waveform_sig_rx =-894;
6579: waveform_sig_rx =-517;
6580: waveform_sig_rx =-806;
6581: waveform_sig_rx =-647;
6582: waveform_sig_rx =-674;
6583: waveform_sig_rx =-712;
6584: waveform_sig_rx =-741;
6585: waveform_sig_rx =-769;
6586: waveform_sig_rx =-588;
6587: waveform_sig_rx =-934;
6588: waveform_sig_rx =-640;
6589: waveform_sig_rx =-648;
6590: waveform_sig_rx =-909;
6591: waveform_sig_rx =-657;
6592: waveform_sig_rx =-606;
6593: waveform_sig_rx =-970;
6594: waveform_sig_rx =-736;
6595: waveform_sig_rx =-581;
6596: waveform_sig_rx =-996;
6597: waveform_sig_rx =-771;
6598: waveform_sig_rx =-615;
6599: waveform_sig_rx =-941;
6600: waveform_sig_rx =-895;
6601: waveform_sig_rx =-594;
6602: waveform_sig_rx =-919;
6603: waveform_sig_rx =-871;
6604: waveform_sig_rx =-778;
6605: waveform_sig_rx =-726;
6606: waveform_sig_rx =-969;
6607: waveform_sig_rx =-844;
6608: waveform_sig_rx =-703;
6609: waveform_sig_rx =-960;
6610: waveform_sig_rx =-951;
6611: waveform_sig_rx =-670;
6612: waveform_sig_rx =-898;
6613: waveform_sig_rx =-1030;
6614: waveform_sig_rx =-666;
6615: waveform_sig_rx =-870;
6616: waveform_sig_rx =-1053;
6617: waveform_sig_rx =-743;
6618: waveform_sig_rx =-830;
6619: waveform_sig_rx =-1058;
6620: waveform_sig_rx =-795;
6621: waveform_sig_rx =-1046;
6622: waveform_sig_rx =-812;
6623: waveform_sig_rx =-952;
6624: waveform_sig_rx =-882;
6625: waveform_sig_rx =-948;
6626: waveform_sig_rx =-994;
6627: waveform_sig_rx =-774;
6628: waveform_sig_rx =-1159;
6629: waveform_sig_rx =-879;
6630: waveform_sig_rx =-824;
6631: waveform_sig_rx =-1188;
6632: waveform_sig_rx =-876;
6633: waveform_sig_rx =-788;
6634: waveform_sig_rx =-1255;
6635: waveform_sig_rx =-867;
6636: waveform_sig_rx =-813;
6637: waveform_sig_rx =-1238;
6638: waveform_sig_rx =-883;
6639: waveform_sig_rx =-879;
6640: waveform_sig_rx =-1126;
6641: waveform_sig_rx =-1048;
6642: waveform_sig_rx =-868;
6643: waveform_sig_rx =-1048;
6644: waveform_sig_rx =-1080;
6645: waveform_sig_rx =-993;
6646: waveform_sig_rx =-878;
6647: waveform_sig_rx =-1191;
6648: waveform_sig_rx =-1001;
6649: waveform_sig_rx =-876;
6650: waveform_sig_rx =-1179;
6651: waveform_sig_rx =-1092;
6652: waveform_sig_rx =-829;
6653: waveform_sig_rx =-1139;
6654: waveform_sig_rx =-1184;
6655: waveform_sig_rx =-836;
6656: waveform_sig_rx =-1134;
6657: waveform_sig_rx =-1163;
6658: waveform_sig_rx =-963;
6659: waveform_sig_rx =-1019;
6660: waveform_sig_rx =-1147;
6661: waveform_sig_rx =-1038;
6662: waveform_sig_rx =-1145;
6663: waveform_sig_rx =-974;
6664: waveform_sig_rx =-1187;
6665: waveform_sig_rx =-980;
6666: waveform_sig_rx =-1163;
6667: waveform_sig_rx =-1148;
6668: waveform_sig_rx =-908;
6669: waveform_sig_rx =-1366;
6670: waveform_sig_rx =-964;
6671: waveform_sig_rx =-992;
6672: waveform_sig_rx =-1358;
6673: waveform_sig_rx =-917;
6674: waveform_sig_rx =-1006;
6675: waveform_sig_rx =-1380;
6676: waveform_sig_rx =-944;
6677: waveform_sig_rx =-1032;
6678: waveform_sig_rx =-1326;
6679: waveform_sig_rx =-986;
6680: waveform_sig_rx =-1051;
6681: waveform_sig_rx =-1198;
6682: waveform_sig_rx =-1187;
6683: waveform_sig_rx =-978;
6684: waveform_sig_rx =-1137;
6685: waveform_sig_rx =-1235;
6686: waveform_sig_rx =-1061;
6687: waveform_sig_rx =-988;
6688: waveform_sig_rx =-1340;
6689: waveform_sig_rx =-1052;
6690: waveform_sig_rx =-1014;
6691: waveform_sig_rx =-1295;
6692: waveform_sig_rx =-1163;
6693: waveform_sig_rx =-979;
6694: waveform_sig_rx =-1257;
6695: waveform_sig_rx =-1228;
6696: waveform_sig_rx =-995;
6697: waveform_sig_rx =-1181;
6698: waveform_sig_rx =-1230;
6699: waveform_sig_rx =-1111;
6700: waveform_sig_rx =-1028;
6701: waveform_sig_rx =-1268;
6702: waveform_sig_rx =-1137;
6703: waveform_sig_rx =-1151;
6704: waveform_sig_rx =-1141;
6705: waveform_sig_rx =-1224;
6706: waveform_sig_rx =-1015;
6707: waveform_sig_rx =-1342;
6708: waveform_sig_rx =-1088;
6709: waveform_sig_rx =-1013;
6710: waveform_sig_rx =-1437;
6711: waveform_sig_rx =-948;
6712: waveform_sig_rx =-1135;
6713: waveform_sig_rx =-1364;
6714: waveform_sig_rx =-974;
6715: waveform_sig_rx =-1125;
6716: waveform_sig_rx =-1388;
6717: waveform_sig_rx =-1002;
6718: waveform_sig_rx =-1099;
6719: waveform_sig_rx =-1355;
6720: waveform_sig_rx =-1061;
6721: waveform_sig_rx =-1099;
6722: waveform_sig_rx =-1246;
6723: waveform_sig_rx =-1250;
6724: waveform_sig_rx =-1016;
6725: waveform_sig_rx =-1189;
6726: waveform_sig_rx =-1308;
6727: waveform_sig_rx =-1056;
6728: waveform_sig_rx =-1057;
6729: waveform_sig_rx =-1409;
6730: waveform_sig_rx =-994;
6731: waveform_sig_rx =-1103;
6732: waveform_sig_rx =-1302;
6733: waveform_sig_rx =-1125;
6734: waveform_sig_rx =-1050;
6735: waveform_sig_rx =-1219;
6736: waveform_sig_rx =-1268;
6737: waveform_sig_rx =-1031;
6738: waveform_sig_rx =-1135;
6739: waveform_sig_rx =-1296;
6740: waveform_sig_rx =-1061;
6741: waveform_sig_rx =-1036;
6742: waveform_sig_rx =-1329;
6743: waveform_sig_rx =-1035;
6744: waveform_sig_rx =-1211;
6745: waveform_sig_rx =-1121;
6746: waveform_sig_rx =-1157;
6747: waveform_sig_rx =-1072;
6748: waveform_sig_rx =-1290;
6749: waveform_sig_rx =-1037;
6750: waveform_sig_rx =-1061;
6751: waveform_sig_rx =-1360;
6752: waveform_sig_rx =-940;
6753: waveform_sig_rx =-1137;
6754: waveform_sig_rx =-1306;
6755: waveform_sig_rx =-953;
6756: waveform_sig_rx =-1112;
6757: waveform_sig_rx =-1323;
6758: waveform_sig_rx =-971;
6759: waveform_sig_rx =-1089;
6760: waveform_sig_rx =-1269;
6761: waveform_sig_rx =-1072;
6762: waveform_sig_rx =-1023;
6763: waveform_sig_rx =-1187;
6764: waveform_sig_rx =-1223;
6765: waveform_sig_rx =-889;
6766: waveform_sig_rx =-1195;
6767: waveform_sig_rx =-1228;
6768: waveform_sig_rx =-936;
6769: waveform_sig_rx =-1090;
6770: waveform_sig_rx =-1250;
6771: waveform_sig_rx =-968;
6772: waveform_sig_rx =-1084;
6773: waveform_sig_rx =-1159;
6774: waveform_sig_rx =-1121;
6775: waveform_sig_rx =-936;
6776: waveform_sig_rx =-1140;
6777: waveform_sig_rx =-1230;
6778: waveform_sig_rx =-883;
6779: waveform_sig_rx =-1130;
6780: waveform_sig_rx =-1229;
6781: waveform_sig_rx =-951;
6782: waveform_sig_rx =-1024;
6783: waveform_sig_rx =-1243;
6784: waveform_sig_rx =-949;
6785: waveform_sig_rx =-1168;
6786: waveform_sig_rx =-1005;
6787: waveform_sig_rx =-1064;
6788: waveform_sig_rx =-992;
6789: waveform_sig_rx =-1175;
6790: waveform_sig_rx =-959;
6791: waveform_sig_rx =-987;
6792: waveform_sig_rx =-1232;
6793: waveform_sig_rx =-861;
6794: waveform_sig_rx =-1067;
6795: waveform_sig_rx =-1162;
6796: waveform_sig_rx =-882;
6797: waveform_sig_rx =-974;
6798: waveform_sig_rx =-1207;
6799: waveform_sig_rx =-899;
6800: waveform_sig_rx =-920;
6801: waveform_sig_rx =-1188;
6802: waveform_sig_rx =-938;
6803: waveform_sig_rx =-857;
6804: waveform_sig_rx =-1162;
6805: waveform_sig_rx =-1025;
6806: waveform_sig_rx =-782;
6807: waveform_sig_rx =-1117;
6808: waveform_sig_rx =-1019;
6809: waveform_sig_rx =-867;
6810: waveform_sig_rx =-943;
6811: waveform_sig_rx =-1098;
6812: waveform_sig_rx =-885;
6813: waveform_sig_rx =-883;
6814: waveform_sig_rx =-1060;
6815: waveform_sig_rx =-984;
6816: waveform_sig_rx =-757;
6817: waveform_sig_rx =-1044;
6818: waveform_sig_rx =-1048;
6819: waveform_sig_rx =-714;
6820: waveform_sig_rx =-1005;
6821: waveform_sig_rx =-1068;
6822: waveform_sig_rx =-765;
6823: waveform_sig_rx =-894;
6824: waveform_sig_rx =-1036;
6825: waveform_sig_rx =-775;
6826: waveform_sig_rx =-1039;
6827: waveform_sig_rx =-789;
6828: waveform_sig_rx =-948;
6829: waveform_sig_rx =-838;
6830: waveform_sig_rx =-976;
6831: waveform_sig_rx =-831;
6832: waveform_sig_rx =-821;
6833: waveform_sig_rx =-1039;
6834: waveform_sig_rx =-741;
6835: waveform_sig_rx =-829;
6836: waveform_sig_rx =-1045;
6837: waveform_sig_rx =-714;
6838: waveform_sig_rx =-764;
6839: waveform_sig_rx =-1110;
6840: waveform_sig_rx =-637;
6841: waveform_sig_rx =-770;
6842: waveform_sig_rx =-1032;
6843: waveform_sig_rx =-682;
6844: waveform_sig_rx =-756;
6845: waveform_sig_rx =-974;
6846: waveform_sig_rx =-810;
6847: waveform_sig_rx =-649;
6848: waveform_sig_rx =-902;
6849: waveform_sig_rx =-836;
6850: waveform_sig_rx =-702;
6851: waveform_sig_rx =-722;
6852: waveform_sig_rx =-922;
6853: waveform_sig_rx =-690;
6854: waveform_sig_rx =-667;
6855: waveform_sig_rx =-894;
6856: waveform_sig_rx =-776;
6857: waveform_sig_rx =-540;
6858: waveform_sig_rx =-880;
6859: waveform_sig_rx =-817;
6860: waveform_sig_rx =-497;
6861: waveform_sig_rx =-834;
6862: waveform_sig_rx =-794;
6863: waveform_sig_rx =-566;
6864: waveform_sig_rx =-726;
6865: waveform_sig_rx =-766;
6866: waveform_sig_rx =-638;
6867: waveform_sig_rx =-790;
6868: waveform_sig_rx =-550;
6869: waveform_sig_rx =-795;
6870: waveform_sig_rx =-540;
6871: waveform_sig_rx =-795;
6872: waveform_sig_rx =-595;
6873: waveform_sig_rx =-543;
6874: waveform_sig_rx =-872;
6875: waveform_sig_rx =-436;
6876: waveform_sig_rx =-620;
6877: waveform_sig_rx =-833;
6878: waveform_sig_rx =-382;
6879: waveform_sig_rx =-610;
6880: waveform_sig_rx =-831;
6881: waveform_sig_rx =-399;
6882: waveform_sig_rx =-587;
6883: waveform_sig_rx =-762;
6884: waveform_sig_rx =-471;
6885: waveform_sig_rx =-523;
6886: waveform_sig_rx =-730;
6887: waveform_sig_rx =-555;
6888: waveform_sig_rx =-449;
6889: waveform_sig_rx =-646;
6890: waveform_sig_rx =-603;
6891: waveform_sig_rx =-484;
6892: waveform_sig_rx =-440;
6893: waveform_sig_rx =-733;
6894: waveform_sig_rx =-420;
6895: waveform_sig_rx =-400;
6896: waveform_sig_rx =-722;
6897: waveform_sig_rx =-420;
6898: waveform_sig_rx =-347;
6899: waveform_sig_rx =-673;
6900: waveform_sig_rx =-478;
6901: waveform_sig_rx =-348;
6902: waveform_sig_rx =-525;
6903: waveform_sig_rx =-535;
6904: waveform_sig_rx =-336;
6905: waveform_sig_rx =-385;
6906: waveform_sig_rx =-566;
6907: waveform_sig_rx =-356;
6908: waveform_sig_rx =-490;
6909: waveform_sig_rx =-345;
6910: waveform_sig_rx =-481;
6911: waveform_sig_rx =-267;
6912: waveform_sig_rx =-580;
6913: waveform_sig_rx =-263;
6914: waveform_sig_rx =-327;
6915: waveform_sig_rx =-608;
6916: waveform_sig_rx =-135;
6917: waveform_sig_rx =-418;
6918: waveform_sig_rx =-534;
6919: waveform_sig_rx =-102;
6920: waveform_sig_rx =-393;
6921: waveform_sig_rx =-524;
6922: waveform_sig_rx =-120;
6923: waveform_sig_rx =-359;
6924: waveform_sig_rx =-443;
6925: waveform_sig_rx =-200;
6926: waveform_sig_rx =-248;
6927: waveform_sig_rx =-436;
6928: waveform_sig_rx =-300;
6929: waveform_sig_rx =-147;
6930: waveform_sig_rx =-339;
6931: waveform_sig_rx =-369;
6932: waveform_sig_rx =-150;
6933: waveform_sig_rx =-181;
6934: waveform_sig_rx =-483;
6935: waveform_sig_rx =-49;
6936: waveform_sig_rx =-207;
6937: waveform_sig_rx =-403;
6938: waveform_sig_rx =-101;
6939: waveform_sig_rx =-142;
6940: waveform_sig_rx =-280;
6941: waveform_sig_rx =-232;
6942: waveform_sig_rx =-58;
6943: waveform_sig_rx =-189;
6944: waveform_sig_rx =-334;
6945: waveform_sig_rx =16;
6946: waveform_sig_rx =-160;
6947: waveform_sig_rx =-290;
6948: waveform_sig_rx =-12;
6949: waveform_sig_rx =-230;
6950: waveform_sig_rx =-54;
6951: waveform_sig_rx =-210;
6952: waveform_sig_rx =1;
6953: waveform_sig_rx =-313;
6954: waveform_sig_rx =49;
6955: waveform_sig_rx =-69;
6956: waveform_sig_rx =-306;
6957: waveform_sig_rx =191;
6958: waveform_sig_rx =-195;
6959: waveform_sig_rx =-212;
6960: waveform_sig_rx =203;
6961: waveform_sig_rx =-165;
6962: waveform_sig_rx =-154;
6963: waveform_sig_rx =122;
6964: waveform_sig_rx =-83;
6965: waveform_sig_rx =-101;
6966: waveform_sig_rx =20;
6967: waveform_sig_rx =98;
6968: waveform_sig_rx =-165;
6969: waveform_sig_rx =-25;
6970: waveform_sig_rx =185;
6971: waveform_sig_rx =-136;
6972: waveform_sig_rx =-35;
6973: waveform_sig_rx =175;
6974: waveform_sig_rx =27;
6975: waveform_sig_rx =-114;
6976: waveform_sig_rx =217;
6977: waveform_sig_rx =79;
6978: waveform_sig_rx =-60;
6979: waveform_sig_rx =153;
6980: waveform_sig_rx =181;
6981: waveform_sig_rx =10;
6982: waveform_sig_rx =34;
6983: waveform_sig_rx =273;
6984: waveform_sig_rx =62;
6985: waveform_sig_rx =-54;
6986: waveform_sig_rx =342;
6987: waveform_sig_rx =129;
6988: waveform_sig_rx =14;
6989: waveform_sig_rx =291;
6990: waveform_sig_rx =39;
6991: waveform_sig_rx =253;
6992: waveform_sig_rx =134;
6993: waveform_sig_rx =271;
6994: waveform_sig_rx =22;
6995: waveform_sig_rx =383;
6996: waveform_sig_rx =155;
6997: waveform_sig_rx =71;
6998: waveform_sig_rx =456;
6999: waveform_sig_rx =78;
7000: waveform_sig_rx =152;
7001: waveform_sig_rx =421;
7002: waveform_sig_rx =182;
7003: waveform_sig_rx =140;
7004: waveform_sig_rx =401;
7005: waveform_sig_rx =281;
7006: waveform_sig_rx =120;
7007: waveform_sig_rx =357;
7008: waveform_sig_rx =421;
7009: waveform_sig_rx =73;
7010: waveform_sig_rx =371;
7011: waveform_sig_rx =458;
7012: waveform_sig_rx =165;
7013: waveform_sig_rx =316;
7014: waveform_sig_rx =434;
7015: waveform_sig_rx =339;
7016: waveform_sig_rx =207;
7017: waveform_sig_rx =498;
7018: waveform_sig_rx =380;
7019: waveform_sig_rx =225;
7020: waveform_sig_rx =416;
7021: waveform_sig_rx =503;
7022: waveform_sig_rx =268;
7023: waveform_sig_rx =339;
7024: waveform_sig_rx =599;
7025: waveform_sig_rx =309;
7026: waveform_sig_rx =284;
7027: waveform_sig_rx =643;
7028: waveform_sig_rx =362;
7029: waveform_sig_rx =343;
7030: waveform_sig_rx =540;
7031: waveform_sig_rx =289;
7032: waveform_sig_rx =589;
7033: waveform_sig_rx =386;
7034: waveform_sig_rx =548;
7035: waveform_sig_rx =337;
7036: waveform_sig_rx =619;
7037: waveform_sig_rx =446;
7038: waveform_sig_rx =364;
7039: waveform_sig_rx =678;
7040: waveform_sig_rx =429;
7041: waveform_sig_rx =398;
7042: waveform_sig_rx =685;
7043: waveform_sig_rx =505;
7044: waveform_sig_rx =329;
7045: waveform_sig_rx =742;
7046: waveform_sig_rx =554;
7047: waveform_sig_rx =358;
7048: waveform_sig_rx =714;
7049: waveform_sig_rx =627;
7050: waveform_sig_rx =340;
7051: waveform_sig_rx =681;
7052: waveform_sig_rx =639;
7053: waveform_sig_rx =467;
7054: waveform_sig_rx =577;
7055: waveform_sig_rx =675;
7056: waveform_sig_rx =626;
7057: waveform_sig_rx =465;
7058: waveform_sig_rx =747;
7059: waveform_sig_rx =683;
7060: waveform_sig_rx =463;
7061: waveform_sig_rx =694;
7062: waveform_sig_rx =809;
7063: waveform_sig_rx =465;
7064: waveform_sig_rx =636;
7065: waveform_sig_rx =848;
7066: waveform_sig_rx =491;
7067: waveform_sig_rx =602;
7068: waveform_sig_rx =841;
7069: waveform_sig_rx =570;
7070: waveform_sig_rx =655;
7071: waveform_sig_rx =718;
7072: waveform_sig_rx =606;
7073: waveform_sig_rx =839;
7074: waveform_sig_rx =591;
7075: waveform_sig_rx =836;
7076: waveform_sig_rx =568;
7077: waveform_sig_rx =874;
7078: waveform_sig_rx =728;
7079: waveform_sig_rx =560;
7080: waveform_sig_rx =942;
7081: waveform_sig_rx =677;
7082: waveform_sig_rx =607;
7083: waveform_sig_rx =1000;
7084: waveform_sig_rx =690;
7085: waveform_sig_rx =577;
7086: waveform_sig_rx =1052;
7087: waveform_sig_rx =699;
7088: waveform_sig_rx =638;
7089: waveform_sig_rx =970;
7090: waveform_sig_rx =801;
7091: waveform_sig_rx =622;
7092: waveform_sig_rx =903;
7093: waveform_sig_rx =858;
7094: waveform_sig_rx =748;
7095: waveform_sig_rx =779;
7096: waveform_sig_rx =949;
7097: waveform_sig_rx =855;
7098: waveform_sig_rx =658;
7099: waveform_sig_rx =1020;
7100: waveform_sig_rx =876;
7101: waveform_sig_rx =666;
7102: waveform_sig_rx =961;
7103: waveform_sig_rx =982;
7104: waveform_sig_rx =672;
7105: waveform_sig_rx =916;
7106: waveform_sig_rx =1021;
7107: waveform_sig_rx =735;
7108: waveform_sig_rx =855;
7109: waveform_sig_rx =1008;
7110: waveform_sig_rx =835;
7111: waveform_sig_rx =863;
7112: waveform_sig_rx =932;
7113: waveform_sig_rx =875;
7114: waveform_sig_rx =990;
7115: waveform_sig_rx =813;
7116: waveform_sig_rx =1066;
7117: waveform_sig_rx =711;
7118: waveform_sig_rx =1115;
7119: waveform_sig_rx =897;
7120: waveform_sig_rx =760;
7121: waveform_sig_rx =1212;
7122: waveform_sig_rx =803;
7123: waveform_sig_rx =823;
7124: waveform_sig_rx =1229;
7125: waveform_sig_rx =781;
7126: waveform_sig_rx =845;
7127: waveform_sig_rx =1206;
7128: waveform_sig_rx =833;
7129: waveform_sig_rx =902;
7130: waveform_sig_rx =1106;
7131: waveform_sig_rx =1002;
7132: waveform_sig_rx =834;
7133: waveform_sig_rx =1035;
7134: waveform_sig_rx =1086;
7135: waveform_sig_rx =898;
7136: waveform_sig_rx =945;
7137: waveform_sig_rx =1156;
7138: waveform_sig_rx =986;
7139: waveform_sig_rx =879;
7140: waveform_sig_rx =1235;
7141: waveform_sig_rx =999;
7142: waveform_sig_rx =846;
7143: waveform_sig_rx =1165;
7144: waveform_sig_rx =1096;
7145: waveform_sig_rx =860;
7146: waveform_sig_rx =1085;
7147: waveform_sig_rx =1119;
7148: waveform_sig_rx =963;
7149: waveform_sig_rx =973;
7150: waveform_sig_rx =1174;
7151: waveform_sig_rx =1046;
7152: waveform_sig_rx =939;
7153: waveform_sig_rx =1151;
7154: waveform_sig_rx =1014;
7155: waveform_sig_rx =1099;
7156: waveform_sig_rx =1071;
7157: waveform_sig_rx =1140;
7158: waveform_sig_rx =876;
7159: waveform_sig_rx =1341;
7160: waveform_sig_rx =944;
7161: waveform_sig_rx =996;
7162: waveform_sig_rx =1334;
7163: waveform_sig_rx =893;
7164: waveform_sig_rx =1063;
7165: waveform_sig_rx =1284;
7166: waveform_sig_rx =957;
7167: waveform_sig_rx =1000;
7168: waveform_sig_rx =1296;
7169: waveform_sig_rx =983;
7170: waveform_sig_rx =1047;
7171: waveform_sig_rx =1224;
7172: waveform_sig_rx =1131;
7173: waveform_sig_rx =941;
7174: waveform_sig_rx =1171;
7175: waveform_sig_rx =1226;
7176: waveform_sig_rx =984;
7177: waveform_sig_rx =1052;
7178: waveform_sig_rx =1314;
7179: waveform_sig_rx =1012;
7180: waveform_sig_rx =1010;
7181: waveform_sig_rx =1325;
7182: waveform_sig_rx =1047;
7183: waveform_sig_rx =1022;
7184: waveform_sig_rx =1224;
7185: waveform_sig_rx =1178;
7186: waveform_sig_rx =1006;
7187: waveform_sig_rx =1125;
7188: waveform_sig_rx =1266;
7189: waveform_sig_rx =1034;
7190: waveform_sig_rx =1023;
7191: waveform_sig_rx =1359;
7192: waveform_sig_rx =1082;
7193: waveform_sig_rx =1048;
7194: waveform_sig_rx =1244;
7195: waveform_sig_rx =1025;
7196: waveform_sig_rx =1218;
7197: waveform_sig_rx =1150;
7198: waveform_sig_rx =1144;
7199: waveform_sig_rx =1011;
7200: waveform_sig_rx =1358;
7201: waveform_sig_rx =992;
7202: waveform_sig_rx =1124;
7203: waveform_sig_rx =1332;
7204: waveform_sig_rx =1004;
7205: waveform_sig_rx =1101;
7206: waveform_sig_rx =1343;
7207: waveform_sig_rx =1032;
7208: waveform_sig_rx =1073;
7209: waveform_sig_rx =1385;
7210: waveform_sig_rx =1015;
7211: waveform_sig_rx =1105;
7212: waveform_sig_rx =1251;
7213: waveform_sig_rx =1187;
7214: waveform_sig_rx =969;
7215: waveform_sig_rx =1219;
7216: waveform_sig_rx =1296;
7217: waveform_sig_rx =975;
7218: waveform_sig_rx =1180;
7219: waveform_sig_rx =1328;
7220: waveform_sig_rx =995;
7221: waveform_sig_rx =1143;
7222: waveform_sig_rx =1261;
7223: waveform_sig_rx =1114;
7224: waveform_sig_rx =1086;
7225: waveform_sig_rx =1176;
7226: waveform_sig_rx =1309;
7227: waveform_sig_rx =956;
7228: waveform_sig_rx =1163;
7229: waveform_sig_rx =1320;
7230: waveform_sig_rx =948;
7231: waveform_sig_rx =1140;
7232: waveform_sig_rx =1325;
7233: waveform_sig_rx =1016;
7234: waveform_sig_rx =1146;
7235: waveform_sig_rx =1197;
7236: waveform_sig_rx =1064;
7237: waveform_sig_rx =1229;
7238: waveform_sig_rx =1082;
7239: waveform_sig_rx =1184;
7240: waveform_sig_rx =1021;
7241: waveform_sig_rx =1332;
7242: waveform_sig_rx =997;
7243: waveform_sig_rx =1121;
7244: waveform_sig_rx =1291;
7245: waveform_sig_rx =1003;
7246: waveform_sig_rx =1103;
7247: waveform_sig_rx =1295;
7248: waveform_sig_rx =1031;
7249: waveform_sig_rx =1016;
7250: waveform_sig_rx =1377;
7251: waveform_sig_rx =1032;
7252: waveform_sig_rx =1024;
7253: waveform_sig_rx =1310;
7254: waveform_sig_rx =1131;
7255: waveform_sig_rx =896;
7256: waveform_sig_rx =1294;
7257: waveform_sig_rx =1144;
7258: waveform_sig_rx =966;
7259: waveform_sig_rx =1161;
7260: waveform_sig_rx =1184;
7261: waveform_sig_rx =1045;
7262: waveform_sig_rx =1058;
7263: waveform_sig_rx =1213;
7264: waveform_sig_rx =1132;
7265: waveform_sig_rx =942;
7266: waveform_sig_rx =1205;
7267: waveform_sig_rx =1212;
7268: waveform_sig_rx =850;
7269: waveform_sig_rx =1210;
7270: waveform_sig_rx =1217;
7271: waveform_sig_rx =906;
7272: waveform_sig_rx =1110;
7273: waveform_sig_rx =1239;
7274: waveform_sig_rx =961;
7275: waveform_sig_rx =1106;
7276: waveform_sig_rx =1080;
7277: waveform_sig_rx =1022;
7278: waveform_sig_rx =1155;
7279: waveform_sig_rx =1015;
7280: waveform_sig_rx =1121;
7281: waveform_sig_rx =935;
7282: waveform_sig_rx =1248;
7283: waveform_sig_rx =948;
7284: waveform_sig_rx =1010;
7285: waveform_sig_rx =1219;
7286: waveform_sig_rx =916;
7287: waveform_sig_rx =986;
7288: waveform_sig_rx =1274;
7289: waveform_sig_rx =884;
7290: waveform_sig_rx =917;
7291: waveform_sig_rx =1325;
7292: waveform_sig_rx =856;
7293: waveform_sig_rx =950;
7294: waveform_sig_rx =1210;
7295: waveform_sig_rx =951;
7296: waveform_sig_rx =870;
7297: waveform_sig_rx =1188;
7298: waveform_sig_rx =996;
7299: waveform_sig_rx =937;
7300: waveform_sig_rx =999;
7301: waveform_sig_rx =1123;
7302: waveform_sig_rx =944;
7303: waveform_sig_rx =893;
7304: waveform_sig_rx =1170;
7305: waveform_sig_rx =962;
7306: waveform_sig_rx =827;
7307: waveform_sig_rx =1137;
7308: waveform_sig_rx =1049;
7309: waveform_sig_rx =757;
7310: waveform_sig_rx =1086;
7311: waveform_sig_rx =1054;
7312: waveform_sig_rx =802;
7313: waveform_sig_rx =987;
7314: waveform_sig_rx =1069;
7315: waveform_sig_rx =822;
7316: waveform_sig_rx =974;
7317: waveform_sig_rx =891;
7318: waveform_sig_rx =933;
7319: waveform_sig_rx =971;
7320: waveform_sig_rx =869;
7321: waveform_sig_rx =1019;
7322: waveform_sig_rx =731;
7323: waveform_sig_rx =1129;
7324: waveform_sig_rx =785;
7325: waveform_sig_rx =834;
7326: waveform_sig_rx =1128;
7327: waveform_sig_rx =687;
7328: waveform_sig_rx =863;
7329: waveform_sig_rx =1138;
7330: waveform_sig_rx =644;
7331: waveform_sig_rx =850;
7332: waveform_sig_rx =1101;
7333: waveform_sig_rx =664;
7334: waveform_sig_rx =847;
7335: waveform_sig_rx =1004;
7336: waveform_sig_rx =807;
7337: waveform_sig_rx =705;
7338: waveform_sig_rx =964;
7339: waveform_sig_rx =850;
7340: waveform_sig_rx =765;
7341: waveform_sig_rx =796;
7342: waveform_sig_rx =976;
7343: waveform_sig_rx =758;
7344: waveform_sig_rx =706;
7345: waveform_sig_rx =1039;
7346: waveform_sig_rx =734;
7347: waveform_sig_rx =655;
7348: waveform_sig_rx =999;
7349: waveform_sig_rx =761;
7350: waveform_sig_rx =631;
7351: waveform_sig_rx =916;
7352: waveform_sig_rx =820;
7353: waveform_sig_rx =666;
7354: waveform_sig_rx =732;
7355: waveform_sig_rx =884;
7356: waveform_sig_rx =669;
7357: waveform_sig_rx =721;
7358: waveform_sig_rx =755;
7359: waveform_sig_rx =741;
7360: waveform_sig_rx =737;
7361: waveform_sig_rx =719;
7362: waveform_sig_rx =742;
7363: waveform_sig_rx =543;
7364: waveform_sig_rx =969;
7365: waveform_sig_rx =507;
7366: waveform_sig_rx =686;
7367: waveform_sig_rx =911;
7368: waveform_sig_rx =440;
7369: waveform_sig_rx =719;
7370: waveform_sig_rx =881;
7371: waveform_sig_rx =422;
7372: waveform_sig_rx =677;
7373: waveform_sig_rx =853;
7374: waveform_sig_rx =450;
7375: waveform_sig_rx =673;
7376: waveform_sig_rx =737;
7377: waveform_sig_rx =601;
7378: waveform_sig_rx =502;
7379: waveform_sig_rx =722;
7380: waveform_sig_rx =649;
7381: waveform_sig_rx =494;
7382: waveform_sig_rx =559;
7383: waveform_sig_rx =785;
7384: waveform_sig_rx =415;
7385: waveform_sig_rx =514;
7386: waveform_sig_rx =766;
7387: waveform_sig_rx =418;
7388: waveform_sig_rx =503;
7389: waveform_sig_rx =682;
7390: waveform_sig_rx =508;
7391: waveform_sig_rx =432;
7392: waveform_sig_rx =594;
7393: waveform_sig_rx =608;
7394: waveform_sig_rx =397;
7395: waveform_sig_rx =471;
7396: waveform_sig_rx =691;
7397: waveform_sig_rx =366;
7398: waveform_sig_rx =500;
7399: waveform_sig_rx =510;
7400: waveform_sig_rx =456;
7401: waveform_sig_rx =487;
7402: waveform_sig_rx =496;
7403: waveform_sig_rx =470;
7404: waveform_sig_rx =336;
7405: waveform_sig_rx =703;
7406: waveform_sig_rx =177;
7407: waveform_sig_rx =478;
7408: waveform_sig_rx =612;
7409: waveform_sig_rx =147;
7410: waveform_sig_rx =533;
7411: waveform_sig_rx =530;
7412: waveform_sig_rx =183;
7413: waveform_sig_rx =430;
7414: waveform_sig_rx =513;
7415: waveform_sig_rx =247;
7416: waveform_sig_rx =346;
7417: waveform_sig_rx =460;
7418: waveform_sig_rx =371;
7419: waveform_sig_rx =143;
7420: waveform_sig_rx =507;
7421: waveform_sig_rx =383;
7422: waveform_sig_rx =189;
7423: waveform_sig_rx =375;
7424: waveform_sig_rx =471;
7425: waveform_sig_rx =144;
7426: waveform_sig_rx =317;
7427: waveform_sig_rx =464;
7428: waveform_sig_rx =164;
7429: waveform_sig_rx =241;
7430: waveform_sig_rx =369;
7431: waveform_sig_rx =297;
7432: waveform_sig_rx =140;
7433: waveform_sig_rx =301;
7434: waveform_sig_rx =360;
7435: waveform_sig_rx =66;
7436: waveform_sig_rx =201;
7437: waveform_sig_rx =417;
7438: waveform_sig_rx =20;
7439: waveform_sig_rx =270;
7440: waveform_sig_rx =188;
7441: waveform_sig_rx =123;
7442: waveform_sig_rx =213;
7443: waveform_sig_rx =183;
7444: waveform_sig_rx =124;
7445: waveform_sig_rx =91;
7446: waveform_sig_rx =365;
7447: waveform_sig_rx =-113;
7448: waveform_sig_rx =248;
7449: waveform_sig_rx =229;
7450: waveform_sig_rx =-78;
7451: waveform_sig_rx =216;
7452: waveform_sig_rx =211;
7453: waveform_sig_rx =-23;
7454: waveform_sig_rx =82;
7455: waveform_sig_rx =255;
7456: waveform_sig_rx =-40;
7457: waveform_sig_rx =3;
7458: waveform_sig_rx =251;
7459: waveform_sig_rx =5;
7460: waveform_sig_rx =-151;
7461: waveform_sig_rx =268;
7462: waveform_sig_rx =-10;
7463: waveform_sig_rx =-79;
7464: waveform_sig_rx =68;
7465: waveform_sig_rx =128;
7466: waveform_sig_rx =-144;
7467: waveform_sig_rx =-10;
7468: waveform_sig_rx =133;
7469: waveform_sig_rx =-117;
7470: waveform_sig_rx =-76;
7471: waveform_sig_rx =60;
7472: waveform_sig_rx =9;
7473: waveform_sig_rx =-211;
7474: waveform_sig_rx =12;
7475: waveform_sig_rx =79;
7476: waveform_sig_rx =-292;
7477: waveform_sig_rx =-16;
7478: waveform_sig_rx =93;
7479: waveform_sig_rx =-334;
7480: waveform_sig_rx =41;
7481: waveform_sig_rx =-204;
7482: waveform_sig_rx =-118;
7483: waveform_sig_rx =-55;
7484: waveform_sig_rx =-178;
7485: waveform_sig_rx =-125;
7486: waveform_sig_rx =-235;
7487: waveform_sig_rx =10;
7488: waveform_sig_rx =-337;
7489: waveform_sig_rx =-103;
7490: waveform_sig_rx =-45;
7491: waveform_sig_rx =-353;
7492: waveform_sig_rx =-128;
7493: waveform_sig_rx =-35;
7494: waveform_sig_rx =-387;
7495: waveform_sig_rx =-227;
7496: waveform_sig_rx =-18;
7497: waveform_sig_rx =-394;
7498: waveform_sig_rx =-272;
7499: waveform_sig_rx =-31;
7500: waveform_sig_rx =-353;
7501: waveform_sig_rx =-397;
7502: waveform_sig_rx =-29;
7503: waveform_sig_rx =-356;
7504: waveform_sig_rx =-342;
7505: waveform_sig_rx =-266;
7506: waveform_sig_rx =-194;
7507: waveform_sig_rx =-428;
7508: waveform_sig_rx =-367;
7509: waveform_sig_rx =-161;
7510: waveform_sig_rx =-419;
7511: waveform_sig_rx =-445;
7512: waveform_sig_rx =-172;
7513: waveform_sig_rx =-341;
7514: waveform_sig_rx =-553;
7515: waveform_sig_rx =-212;
7516: waveform_sig_rx =-308;
7517: waveform_sig_rx =-580;
7518: waveform_sig_rx =-279;
7519: waveform_sig_rx =-302;
7520: waveform_sig_rx =-569;
7521: waveform_sig_rx =-273;
7522: waveform_sig_rx =-507;
7523: waveform_sig_rx =-350;
7524: waveform_sig_rx =-417;
7525: waveform_sig_rx =-441;
7526: waveform_sig_rx =-389;
7527: waveform_sig_rx =-566;
7528: waveform_sig_rx =-234;
7529: waveform_sig_rx =-634;
7530: waveform_sig_rx =-438;
7531: waveform_sig_rx =-298;
7532: waveform_sig_rx =-691;
7533: waveform_sig_rx =-431;
7534: waveform_sig_rx =-308;
7535: waveform_sig_rx =-730;
7536: waveform_sig_rx =-472;
7537: waveform_sig_rx =-300;
7538: waveform_sig_rx =-738;
7539: waveform_sig_rx =-506;
7540: waveform_sig_rx =-363;
7541: waveform_sig_rx =-669;
7542: waveform_sig_rx =-624;
7543: waveform_sig_rx =-375;
7544: waveform_sig_rx =-629;
7545: waveform_sig_rx =-612;
7546: waveform_sig_rx =-578;
7547: waveform_sig_rx =-425;
7548: waveform_sig_rx =-718;
7549: waveform_sig_rx =-620;
7550: waveform_sig_rx =-388;
7551: waveform_sig_rx =-732;
7552: waveform_sig_rx =-718;
7553: waveform_sig_rx =-411;
7554: waveform_sig_rx =-670;
7555: waveform_sig_rx =-784;
7556: waveform_sig_rx =-454;
7557: waveform_sig_rx =-646;
7558: waveform_sig_rx =-769;
7559: waveform_sig_rx =-589;
7560: waveform_sig_rx =-565;
7561: waveform_sig_rx =-784;
7562: waveform_sig_rx =-628;
7563: waveform_sig_rx =-752;
7564: waveform_sig_rx =-633;
7565: waveform_sig_rx =-753;
7566: waveform_sig_rx =-659;
7567: waveform_sig_rx =-725;
7568: waveform_sig_rx =-827;
7569: waveform_sig_rx =-494;
7570: waveform_sig_rx =-966;
7571: waveform_sig_rx =-674;
7572: waveform_sig_rx =-572;
7573: waveform_sig_rx =-1011;
7574: waveform_sig_rx =-651;
7575: waveform_sig_rx =-591;
7576: waveform_sig_rx =-1053;
7577: waveform_sig_rx =-664;
7578: waveform_sig_rx =-631;
7579: waveform_sig_rx =-1006;
7580: waveform_sig_rx =-689;
7581: waveform_sig_rx =-705;
7582: waveform_sig_rx =-870;
7583: waveform_sig_rx =-899;
7584: waveform_sig_rx =-686;
7585: waveform_sig_rx =-819;
7586: waveform_sig_rx =-909;
7587: waveform_sig_rx =-807;
7588: waveform_sig_rx =-663;
7589: waveform_sig_rx =-1027;
7590: waveform_sig_rx =-823;
7591: waveform_sig_rx =-667;
7592: waveform_sig_rx =-1011;
7593: waveform_sig_rx =-909;
7594: waveform_sig_rx =-674;
7595: waveform_sig_rx =-944;
7596: waveform_sig_rx =-979;
7597: waveform_sig_rx =-728;
7598: waveform_sig_rx =-893;
7599: waveform_sig_rx =-964;
7600: waveform_sig_rx =-881;
7601: waveform_sig_rx =-758;
7602: waveform_sig_rx =-1016;
7603: waveform_sig_rx =-896;
7604: waveform_sig_rx =-880;
7605: waveform_sig_rx =-907;
7606: waveform_sig_rx =-968;
7607: waveform_sig_rx =-820;
7608: waveform_sig_rx =-1037;
7609: waveform_sig_rx =-952;
7610: waveform_sig_rx =-744;
7611: waveform_sig_rx =-1236;
7612: waveform_sig_rx =-783;
7613: waveform_sig_rx =-877;
7614: waveform_sig_rx =-1195;
7615: waveform_sig_rx =-819;
7616: waveform_sig_rx =-874;
7617: waveform_sig_rx =-1193;
7618: waveform_sig_rx =-869;
7619: waveform_sig_rx =-859;
7620: waveform_sig_rx =-1185;
7621: waveform_sig_rx =-931;
7622: waveform_sig_rx =-911;
7623: waveform_sig_rx =-1061;
7624: waveform_sig_rx =-1131;
7625: waveform_sig_rx =-852;
7626: waveform_sig_rx =-1004;
7627: waveform_sig_rx =-1163;
7628: waveform_sig_rx =-967;
7629: waveform_sig_rx =-869;
7630: waveform_sig_rx =-1247;
7631: waveform_sig_rx =-929;
7632: waveform_sig_rx =-907;
7633: waveform_sig_rx =-1204;
7634: waveform_sig_rx =-1022;
7635: waveform_sig_rx =-939;
7636: waveform_sig_rx =-1069;
7637: waveform_sig_rx =-1152;
7638: waveform_sig_rx =-958;
7639: waveform_sig_rx =-971;
7640: waveform_sig_rx =-1231;
7641: waveform_sig_rx =-1024;
7642: waveform_sig_rx =-889;
7643: waveform_sig_rx =-1283;
7644: waveform_sig_rx =-959;
7645: waveform_sig_rx =-1107;
7646: waveform_sig_rx =-1089;
7647: waveform_sig_rx =-1053;
7648: waveform_sig_rx =-1034;
7649: waveform_sig_rx =-1192;
7650: waveform_sig_rx =-1038;
7651: waveform_sig_rx =-965;
7652: waveform_sig_rx =-1326;
7653: waveform_sig_rx =-925;
7654: waveform_sig_rx =-1049;
7655: waveform_sig_rx =-1279;
7656: waveform_sig_rx =-959;
7657: waveform_sig_rx =-1016;
7658: waveform_sig_rx =-1326;
7659: waveform_sig_rx =-1008;
7660: waveform_sig_rx =-1019;
7661: waveform_sig_rx =-1301;
7662: waveform_sig_rx =-1078;
7663: waveform_sig_rx =-1023;
7664: waveform_sig_rx =-1166;
7665: waveform_sig_rx =-1279;
7666: waveform_sig_rx =-907;
7667: waveform_sig_rx =-1165;
7668: waveform_sig_rx =-1292;
7669: waveform_sig_rx =-989;
7670: waveform_sig_rx =-1078;
7671: waveform_sig_rx =-1306;
7672: waveform_sig_rx =-1023;
7673: waveform_sig_rx =-1108;
7674: waveform_sig_rx =-1202;
7675: waveform_sig_rx =-1198;
7676: waveform_sig_rx =-1011;
7677: waveform_sig_rx =-1123;
7678: waveform_sig_rx =-1325;
7679: waveform_sig_rx =-972;
7680: waveform_sig_rx =-1119;
7681: waveform_sig_rx =-1339;
7682: waveform_sig_rx =-1018;
7683: waveform_sig_rx =-1054;
7684: waveform_sig_rx =-1332;
7685: waveform_sig_rx =-1028;
7686: waveform_sig_rx =-1262;
7687: waveform_sig_rx =-1110;
7688: waveform_sig_rx =-1154;
7689: waveform_sig_rx =-1124;
7690: waveform_sig_rx =-1220;
7691: waveform_sig_rx =-1139;
7692: waveform_sig_rx =-1044;
7693: waveform_sig_rx =-1363;
7694: waveform_sig_rx =-1010;
7695: waveform_sig_rx =-1131;
7696: waveform_sig_rx =-1329;
7697: waveform_sig_rx =-1040;
7698: waveform_sig_rx =-1065;
7699: waveform_sig_rx =-1335;
7700: waveform_sig_rx =-1091;
7701: waveform_sig_rx =-1028;
7702: waveform_sig_rx =-1344;
7703: waveform_sig_rx =-1118;
7704: waveform_sig_rx =-988;
7705: waveform_sig_rx =-1308;
7706: waveform_sig_rx =-1269;
7707: waveform_sig_rx =-933;
7708: waveform_sig_rx =-1304;
7709: waveform_sig_rx =-1211;
7710: waveform_sig_rx =-1086;
7711: waveform_sig_rx =-1138;
7712: waveform_sig_rx =-1250;
7713: waveform_sig_rx =-1151;
7714: waveform_sig_rx =-1041;
7715: waveform_sig_rx =-1233;
7716: waveform_sig_rx =-1256;
7717: waveform_sig_rx =-939;
7718: waveform_sig_rx =-1252;
7719: waveform_sig_rx =-1277;
7720: waveform_sig_rx =-948;
7721: waveform_sig_rx =-1197;
7722: waveform_sig_rx =-1280;
7723: waveform_sig_rx =-1044;
7724: waveform_sig_rx =-1073;
7725: waveform_sig_rx =-1308;
7726: waveform_sig_rx =-1033;
7727: waveform_sig_rx =-1234;
7728: waveform_sig_rx =-1088;
7729: waveform_sig_rx =-1149;
7730: waveform_sig_rx =-1118;
7731: waveform_sig_rx =-1229;
7732: waveform_sig_rx =-1116;
7733: waveform_sig_rx =-1054;
7734: waveform_sig_rx =-1322;
7735: waveform_sig_rx =-1037;
7736: waveform_sig_rx =-1085;
7737: waveform_sig_rx =-1302;
7738: waveform_sig_rx =-1043;
7739: waveform_sig_rx =-974;
7740: waveform_sig_rx =-1407;
7741: waveform_sig_rx =-986;
7742: waveform_sig_rx =-995;
7743: waveform_sig_rx =-1386;
7744: waveform_sig_rx =-961;
7745: waveform_sig_rx =-1026;
7746: waveform_sig_rx =-1257;
7747: waveform_sig_rx =-1138;
7748: waveform_sig_rx =-969;
7749: waveform_sig_rx =-1178;
7750: waveform_sig_rx =-1178;
7751: waveform_sig_rx =-1057;
7752: waveform_sig_rx =-996;
7753: waveform_sig_rx =-1272;
7754: waveform_sig_rx =-1062;
7755: waveform_sig_rx =-969;
7756: waveform_sig_rx =-1234;
7757: waveform_sig_rx =-1136;
7758: waveform_sig_rx =-872;
7759: waveform_sig_rx =-1211;
7760: waveform_sig_rx =-1192;
7761: waveform_sig_rx =-883;
7762: waveform_sig_rx =-1148;
7763: waveform_sig_rx =-1174;
7764: waveform_sig_rx =-962;
7765: waveform_sig_rx =-1028;
7766: waveform_sig_rx =-1178;
7767: waveform_sig_rx =-973;
7768: waveform_sig_rx =-1168;
7769: waveform_sig_rx =-947;
7770: waveform_sig_rx =-1133;
7771: waveform_sig_rx =-970;
7772: waveform_sig_rx =-1114;
7773: waveform_sig_rx =-1059;
7774: waveform_sig_rx =-913;
7775: waveform_sig_rx =-1279;
7776: waveform_sig_rx =-905;
7777: waveform_sig_rx =-945;
7778: waveform_sig_rx =-1273;
7779: waveform_sig_rx =-832;
7780: waveform_sig_rx =-944;
7781: waveform_sig_rx =-1301;
7782: waveform_sig_rx =-782;
7783: waveform_sig_rx =-963;
7784: waveform_sig_rx =-1206;
7785: waveform_sig_rx =-860;
7786: waveform_sig_rx =-957;
7787: waveform_sig_rx =-1090;
7788: waveform_sig_rx =-1018;
7789: waveform_sig_rx =-840;
7790: waveform_sig_rx =-1026;
7791: waveform_sig_rx =-1065;
7792: waveform_sig_rx =-902;
7793: waveform_sig_rx =-872;
7794: waveform_sig_rx =-1168;
7795: waveform_sig_rx =-866;
7796: waveform_sig_rx =-824;
7797: waveform_sig_rx =-1117;
7798: waveform_sig_rx =-934;
7799: waveform_sig_rx =-758;
7800: waveform_sig_rx =-1076;
7801: waveform_sig_rx =-992;
7802: waveform_sig_rx =-771;
7803: waveform_sig_rx =-987;
7804: waveform_sig_rx =-1005;
7805: waveform_sig_rx =-865;
7806: waveform_sig_rx =-844;
7807: waveform_sig_rx =-1029;
7808: waveform_sig_rx =-850;
7809: waveform_sig_rx =-945;
7810: waveform_sig_rx =-826;
7811: waveform_sig_rx =-978;
7812: waveform_sig_rx =-755;
7813: waveform_sig_rx =-1050;
7814: waveform_sig_rx =-808;
7815: waveform_sig_rx =-742;
7816: waveform_sig_rx =-1145;
7817: waveform_sig_rx =-634;
7818: waveform_sig_rx =-857;
7819: waveform_sig_rx =-1065;
7820: waveform_sig_rx =-614;
7821: waveform_sig_rx =-855;
7822: waveform_sig_rx =-1022;
7823: waveform_sig_rx =-647;
7824: waveform_sig_rx =-810;
7825: waveform_sig_rx =-968;
7826: waveform_sig_rx =-740;
7827: waveform_sig_rx =-760;
7828: waveform_sig_rx =-922;
7829: waveform_sig_rx =-846;
7830: waveform_sig_rx =-638;
7831: waveform_sig_rx =-840;
7832: waveform_sig_rx =-902;
7833: waveform_sig_rx =-697;
7834: waveform_sig_rx =-686;
7835: waveform_sig_rx =-1010;
7836: waveform_sig_rx =-605;
7837: waveform_sig_rx =-674;
7838: waveform_sig_rx =-938;
7839: waveform_sig_rx =-681;
7840: waveform_sig_rx =-662;
7841: waveform_sig_rx =-822;
7842: waveform_sig_rx =-795;
7843: waveform_sig_rx =-617;
7844: waveform_sig_rx =-697;
7845: waveform_sig_rx =-875;
7846: waveform_sig_rx =-588;
7847: waveform_sig_rx =-601;
7848: waveform_sig_rx =-875;
7849: waveform_sig_rx =-552;
7850: waveform_sig_rx =-781;
7851: waveform_sig_rx =-609;
7852: waveform_sig_rx =-710;
7853: waveform_sig_rx =-575;
7854: waveform_sig_rx =-838;
7855: waveform_sig_rx =-545;
7856: waveform_sig_rx =-593;
7857: waveform_sig_rx =-887;
7858: waveform_sig_rx =-392;
7859: waveform_sig_rx =-703;
7860: waveform_sig_rx =-784;
7861: waveform_sig_rx =-405;
7862: waveform_sig_rx =-673;
7863: waveform_sig_rx =-736;
7864: waveform_sig_rx =-454;
7865: waveform_sig_rx =-572;
7866: waveform_sig_rx =-702;
7867: waveform_sig_rx =-543;
7868: waveform_sig_rx =-433;
7869: waveform_sig_rx =-716;
7870: waveform_sig_rx =-626;
7871: waveform_sig_rx =-356;
7872: waveform_sig_rx =-657;
7873: waveform_sig_rx =-612;
7874: waveform_sig_rx =-414;
7875: waveform_sig_rx =-498;
7876: waveform_sig_rx =-702;
7877: waveform_sig_rx =-374;
7878: waveform_sig_rx =-462;
7879: waveform_sig_rx =-652;
7880: waveform_sig_rx =-438;
7881: waveform_sig_rx =-408;
7882: waveform_sig_rx =-531;
7883: waveform_sig_rx =-563;
7884: waveform_sig_rx =-323;
7885: waveform_sig_rx =-451;
7886: waveform_sig_rx =-673;
7887: waveform_sig_rx =-258;
7888: waveform_sig_rx =-408;
7889: waveform_sig_rx =-608;
7890: waveform_sig_rx =-256;
7891: waveform_sig_rx =-564;
7892: waveform_sig_rx =-318;
7893: waveform_sig_rx =-426;
7894: waveform_sig_rx =-349;
7895: waveform_sig_rx =-532;
7896: waveform_sig_rx =-274;
7897: waveform_sig_rx =-381;
7898: waveform_sig_rx =-544;
7899: waveform_sig_rx =-173;
7900: waveform_sig_rx =-437;
7901: waveform_sig_rx =-455;
7902: waveform_sig_rx =-191;
7903: waveform_sig_rx =-373;
7904: waveform_sig_rx =-484;
7905: waveform_sig_rx =-198;
7906: waveform_sig_rx =-263;
7907: waveform_sig_rx =-477;
7908: waveform_sig_rx =-221;
7909: waveform_sig_rx =-157;
7910: waveform_sig_rx =-495;
7911: waveform_sig_rx =-276;
7912: waveform_sig_rx =-118;
7913: waveform_sig_rx =-423;
7914: waveform_sig_rx =-299;
7915: waveform_sig_rx =-173;
7916: waveform_sig_rx =-227;
7917: waveform_sig_rx =-398;
7918: waveform_sig_rx =-120;
7919: waveform_sig_rx =-202;
7920: waveform_sig_rx =-340;
7921: waveform_sig_rx =-204;
7922: waveform_sig_rx =-89;
7923: waveform_sig_rx =-270;
7924: waveform_sig_rx =-322;
7925: waveform_sig_rx =18;
7926: waveform_sig_rx =-249;
7927: waveform_sig_rx =-356;
7928: waveform_sig_rx =63;
7929: waveform_sig_rx =-197;
7930: waveform_sig_rx =-255;
7931: waveform_sig_rx =10;
7932: waveform_sig_rx =-307;
7933: waveform_sig_rx =21;
7934: waveform_sig_rx =-202;
7935: waveform_sig_rx =-56;
7936: waveform_sig_rx =-215;
7937: waveform_sig_rx =-8;
7938: waveform_sig_rx =-68;
7939: waveform_sig_rx =-255;
7940: waveform_sig_rx =96;
7941: waveform_sig_rx =-102;
7942: waveform_sig_rx =-207;
7943: waveform_sig_rx =124;
7944: waveform_sig_rx =-47;
7945: waveform_sig_rx =-251;
7946: waveform_sig_rx =121;
7947: waveform_sig_rx =10;
7948: waveform_sig_rx =-230;
7949: waveform_sig_rx =110;
7950: waveform_sig_rx =103;
7951: waveform_sig_rx =-223;
7952: waveform_sig_rx =63;
7953: waveform_sig_rx =152;
7954: waveform_sig_rx =-110;
7955: waveform_sig_rx =32;
7956: waveform_sig_rx =110;
7957: waveform_sig_rx =88;
7958: waveform_sig_rx =-83;
7959: waveform_sig_rx =163;
7960: waveform_sig_rx =143;
7961: waveform_sig_rx =-79;
7962: waveform_sig_rx =93;
7963: waveform_sig_rx =267;
7964: waveform_sig_rx =-64;
7965: waveform_sig_rx =23;
7966: waveform_sig_rx =325;
7967: waveform_sig_rx =-16;
7968: waveform_sig_rx =32;
7969: waveform_sig_rx =306;
7970: waveform_sig_rx =73;
7971: waveform_sig_rx =80;
7972: waveform_sig_rx =228;
7973: waveform_sig_rx =40;
7974: waveform_sig_rx =306;
7975: waveform_sig_rx =61;
7976: waveform_sig_rx =303;
7977: waveform_sig_rx =50;
7978: waveform_sig_rx =293;
7979: waveform_sig_rx =242;
7980: waveform_sig_rx =24;
7981: waveform_sig_rx =397;
7982: waveform_sig_rx =174;
7983: waveform_sig_rx =48;
7984: waveform_sig_rx =433;
7985: waveform_sig_rx =245;
7986: waveform_sig_rx =9;
7987: waveform_sig_rx =468;
7988: waveform_sig_rx =265;
7989: waveform_sig_rx =50;
7990: waveform_sig_rx =450;
7991: waveform_sig_rx =319;
7992: waveform_sig_rx =91;
7993: waveform_sig_rx =379;
7994: waveform_sig_rx =364;
7995: waveform_sig_rx =244;
7996: waveform_sig_rx =273;
7997: waveform_sig_rx =388;
7998: waveform_sig_rx =414;
7999: waveform_sig_rx =114;
8000: waveform_sig_rx =480;
8001: waveform_sig_rx =413;
8002: waveform_sig_rx =143;
8003: waveform_sig_rx =444;
8004: waveform_sig_rx =493;
8005: waveform_sig_rx =212;
8006: waveform_sig_rx =377;
8007: waveform_sig_rx =555;
8008: waveform_sig_rx =285;
8009: waveform_sig_rx =316;
8010: waveform_sig_rx =542;
8011: waveform_sig_rx =377;
8012: waveform_sig_rx =367;
8013: waveform_sig_rx =469;
8014: waveform_sig_rx =374;
8015: waveform_sig_rx =560;
8016: waveform_sig_rx =344;
8017: waveform_sig_rx =622;
8018: waveform_sig_rx =280;
8019: waveform_sig_rx =608;
8020: waveform_sig_rx =511;
8021: waveform_sig_rx =262;
8022: waveform_sig_rx =730;
8023: waveform_sig_rx =432;
8024: waveform_sig_rx =299;
8025: waveform_sig_rx =776;
8026: waveform_sig_rx =415;
8027: waveform_sig_rx =314;
8028: waveform_sig_rx =769;
8029: waveform_sig_rx =451;
8030: waveform_sig_rx =404;
8031: waveform_sig_rx =671;
8032: waveform_sig_rx =572;
8033: waveform_sig_rx =418;
8034: waveform_sig_rx =593;
8035: waveform_sig_rx =663;
8036: waveform_sig_rx =517;
8037: waveform_sig_rx =494;
8038: waveform_sig_rx =719;
8039: waveform_sig_rx =624;
8040: waveform_sig_rx =405;
8041: waveform_sig_rx =802;
8042: waveform_sig_rx =637;
8043: waveform_sig_rx =424;
8044: waveform_sig_rx =750;
8045: waveform_sig_rx =719;
8046: waveform_sig_rx =470;
8047: waveform_sig_rx =661;
8048: waveform_sig_rx =774;
8049: waveform_sig_rx =587;
8050: waveform_sig_rx =587;
8051: waveform_sig_rx =785;
8052: waveform_sig_rx =675;
8053: waveform_sig_rx =570;
8054: waveform_sig_rx =753;
8055: waveform_sig_rx =662;
8056: waveform_sig_rx =735;
8057: waveform_sig_rx =661;
8058: waveform_sig_rx =841;
8059: waveform_sig_rx =484;
8060: waveform_sig_rx =936;
8061: waveform_sig_rx =686;
8062: waveform_sig_rx =546;
8063: waveform_sig_rx =1018;
8064: waveform_sig_rx =591;
8065: waveform_sig_rx =643;
8066: waveform_sig_rx =980;
8067: waveform_sig_rx =639;
8068: waveform_sig_rx =639;
8069: waveform_sig_rx =959;
8070: waveform_sig_rx =689;
8071: waveform_sig_rx =662;
8072: waveform_sig_rx =883;
8073: waveform_sig_rx =838;
8074: waveform_sig_rx =646;
8075: waveform_sig_rx =802;
8076: waveform_sig_rx =933;
8077: waveform_sig_rx =709;
8078: waveform_sig_rx =723;
8079: waveform_sig_rx =994;
8080: waveform_sig_rx =791;
8081: waveform_sig_rx =667;
8082: waveform_sig_rx =1065;
8083: waveform_sig_rx =808;
8084: waveform_sig_rx =723;
8085: waveform_sig_rx =959;
8086: waveform_sig_rx =946;
8087: waveform_sig_rx =765;
8088: waveform_sig_rx =860;
8089: waveform_sig_rx =1010;
8090: waveform_sig_rx =832;
8091: waveform_sig_rx =752;
8092: waveform_sig_rx =1055;
8093: waveform_sig_rx =884;
8094: waveform_sig_rx =754;
8095: waveform_sig_rx =1045;
8096: waveform_sig_rx =791;
8097: waveform_sig_rx =958;
8098: waveform_sig_rx =906;
8099: waveform_sig_rx =943;
8100: waveform_sig_rx =766;
8101: waveform_sig_rx =1126;
8102: waveform_sig_rx =824;
8103: waveform_sig_rx =845;
8104: waveform_sig_rx =1142;
8105: waveform_sig_rx =813;
8106: waveform_sig_rx =870;
8107: waveform_sig_rx =1142;
8108: waveform_sig_rx =866;
8109: waveform_sig_rx =816;
8110: waveform_sig_rx =1192;
8111: waveform_sig_rx =856;
8112: waveform_sig_rx =887;
8113: waveform_sig_rx =1074;
8114: waveform_sig_rx =1045;
8115: waveform_sig_rx =829;
8116: waveform_sig_rx =985;
8117: waveform_sig_rx =1189;
8118: waveform_sig_rx =823;
8119: waveform_sig_rx =972;
8120: waveform_sig_rx =1219;
8121: waveform_sig_rx =888;
8122: waveform_sig_rx =938;
8123: waveform_sig_rx =1151;
8124: waveform_sig_rx =980;
8125: waveform_sig_rx =942;
8126: waveform_sig_rx =1012;
8127: waveform_sig_rx =1163;
8128: waveform_sig_rx =847;
8129: waveform_sig_rx =989;
8130: waveform_sig_rx =1240;
8131: waveform_sig_rx =875;
8132: waveform_sig_rx =969;
8133: waveform_sig_rx =1227;
8134: waveform_sig_rx =945;
8135: waveform_sig_rx =988;
8136: waveform_sig_rx =1132;
8137: waveform_sig_rx =925;
8138: waveform_sig_rx =1164;
8139: waveform_sig_rx =1014;
8140: waveform_sig_rx =1083;
8141: waveform_sig_rx =939;
8142: waveform_sig_rx =1248;
8143: waveform_sig_rx =958;
8144: waveform_sig_rx =993;
8145: waveform_sig_rx =1236;
8146: waveform_sig_rx =963;
8147: waveform_sig_rx =1023;
8148: waveform_sig_rx =1253;
8149: waveform_sig_rx =1018;
8150: waveform_sig_rx =921;
8151: waveform_sig_rx =1313;
8152: waveform_sig_rx =1033;
8153: waveform_sig_rx =945;
8154: waveform_sig_rx =1239;
8155: waveform_sig_rx =1159;
8156: waveform_sig_rx =878;
8157: waveform_sig_rx =1206;
8158: waveform_sig_rx =1202;
8159: waveform_sig_rx =933;
8160: waveform_sig_rx =1152;
8161: waveform_sig_rx =1197;
8162: waveform_sig_rx =1041;
8163: waveform_sig_rx =1044;
8164: waveform_sig_rx =1192;
8165: waveform_sig_rx =1159;
8166: waveform_sig_rx =954;
8167: waveform_sig_rx =1169;
8168: waveform_sig_rx =1289;
8169: waveform_sig_rx =875;
8170: waveform_sig_rx =1164;
8171: waveform_sig_rx =1275;
8172: waveform_sig_rx =956;
8173: waveform_sig_rx =1092;
8174: waveform_sig_rx =1284;
8175: waveform_sig_rx =1050;
8176: waveform_sig_rx =1077;
8177: waveform_sig_rx =1193;
8178: waveform_sig_rx =1028;
8179: waveform_sig_rx =1236;
8180: waveform_sig_rx =1071;
8181: waveform_sig_rx =1176;
8182: waveform_sig_rx =990;
8183: waveform_sig_rx =1306;
8184: waveform_sig_rx =1068;
8185: waveform_sig_rx =1074;
8186: waveform_sig_rx =1297;
8187: waveform_sig_rx =1073;
8188: waveform_sig_rx =1040;
8189: waveform_sig_rx =1356;
8190: waveform_sig_rx =1075;
8191: waveform_sig_rx =940;
8192: waveform_sig_rx =1444;
8193: waveform_sig_rx =1017;
8194: waveform_sig_rx =1011;
8195: waveform_sig_rx =1371;
8196: waveform_sig_rx =1101;
8197: waveform_sig_rx =995;
8198: waveform_sig_rx =1266;
8199: waveform_sig_rx =1159;
8200: waveform_sig_rx =1078;
8201: waveform_sig_rx =1124;
8202: waveform_sig_rx =1266;
8203: waveform_sig_rx =1136;
8204: waveform_sig_rx =1003;
8205: waveform_sig_rx =1305;
8206: waveform_sig_rx =1140;
8207: waveform_sig_rx =973;
8208: waveform_sig_rx =1269;
8209: waveform_sig_rx =1241;
8210: waveform_sig_rx =945;
8211: waveform_sig_rx =1228;
8212: waveform_sig_rx =1277;
8213: waveform_sig_rx =998;
8214: waveform_sig_rx =1156;
8215: waveform_sig_rx =1293;
8216: waveform_sig_rx =1058;
8217: waveform_sig_rx =1153;
8218: waveform_sig_rx =1167;
8219: waveform_sig_rx =1085;
8220: waveform_sig_rx =1230;
8221: waveform_sig_rx =1037;
8222: waveform_sig_rx =1260;
8223: waveform_sig_rx =941;
8224: waveform_sig_rx =1311;
8225: waveform_sig_rx =1074;
8226: waveform_sig_rx =981;
8227: waveform_sig_rx =1369;
8228: waveform_sig_rx =975;
8229: waveform_sig_rx =1003;
8230: waveform_sig_rx =1425;
8231: waveform_sig_rx =928;
8232: waveform_sig_rx =1031;
8233: waveform_sig_rx =1417;
8234: waveform_sig_rx =935;
8235: waveform_sig_rx =1111;
8236: waveform_sig_rx =1251;
8237: waveform_sig_rx =1109;
8238: waveform_sig_rx =998;
8239: waveform_sig_rx =1199;
8240: waveform_sig_rx =1202;
8241: waveform_sig_rx =1007;
8242: waveform_sig_rx =1064;
8243: waveform_sig_rx =1262;
8244: waveform_sig_rx =1030;
8245: waveform_sig_rx =964;
8246: waveform_sig_rx =1291;
8247: waveform_sig_rx =1077;
8248: waveform_sig_rx =950;
8249: waveform_sig_rx =1263;
8250: waveform_sig_rx =1161;
8251: waveform_sig_rx =902;
8252: waveform_sig_rx =1184;
8253: waveform_sig_rx =1174;
8254: waveform_sig_rx =983;
8255: waveform_sig_rx =1073;
8256: waveform_sig_rx =1222;
8257: waveform_sig_rx =1044;
8258: waveform_sig_rx =1038;
8259: waveform_sig_rx =1110;
8260: waveform_sig_rx =1053;
8261: waveform_sig_rx =1099;
8262: waveform_sig_rx =1050;
8263: waveform_sig_rx =1154;
8264: waveform_sig_rx =869;
8265: waveform_sig_rx =1317;
8266: waveform_sig_rx =900;
8267: waveform_sig_rx =978;
8268: waveform_sig_rx =1328;
8269: waveform_sig_rx =815;
8270: waveform_sig_rx =1031;
8271: waveform_sig_rx =1266;
8272: waveform_sig_rx =819;
8273: waveform_sig_rx =980;
8274: waveform_sig_rx =1245;
8275: waveform_sig_rx =875;
8276: waveform_sig_rx =998;
8277: waveform_sig_rx =1138;
8278: waveform_sig_rx =1024;
8279: waveform_sig_rx =877;
8280: waveform_sig_rx =1107;
8281: waveform_sig_rx =1091;
8282: waveform_sig_rx =904;
8283: waveform_sig_rx =956;
8284: waveform_sig_rx =1178;
8285: waveform_sig_rx =882;
8286: waveform_sig_rx =893;
8287: waveform_sig_rx =1211;
8288: waveform_sig_rx =883;
8289: waveform_sig_rx =888;
8290: waveform_sig_rx =1135;
8291: waveform_sig_rx =975;
8292: waveform_sig_rx =866;
8293: waveform_sig_rx =1023;
8294: waveform_sig_rx =1058;
8295: waveform_sig_rx =879;
8296: waveform_sig_rx =881;
8297: waveform_sig_rx =1161;
8298: waveform_sig_rx =850;
8299: waveform_sig_rx =884;
8300: waveform_sig_rx =1028;
8301: waveform_sig_rx =877;
8302: waveform_sig_rx =978;
8303: waveform_sig_rx =944;
8304: waveform_sig_rx =937;
8305: waveform_sig_rx =772;
8306: waveform_sig_rx =1158;
8307: waveform_sig_rx =698;
8308: waveform_sig_rx =906;
8309: waveform_sig_rx =1079;
8310: waveform_sig_rx =673;
8311: waveform_sig_rx =934;
8312: waveform_sig_rx =1062;
8313: waveform_sig_rx =713;
8314: waveform_sig_rx =844;
8315: waveform_sig_rx =1054;
8316: waveform_sig_rx =739;
8317: waveform_sig_rx =836;
8318: waveform_sig_rx =960;
8319: waveform_sig_rx =895;
8320: waveform_sig_rx =660;
8321: waveform_sig_rx =952;
8322: waveform_sig_rx =917;
8323: waveform_sig_rx =673;
8324: waveform_sig_rx =829;
8325: waveform_sig_rx =993;
8326: waveform_sig_rx =666;
8327: waveform_sig_rx =783;
8328: waveform_sig_rx =988;
8329: waveform_sig_rx =705;
8330: waveform_sig_rx =727;
8331: waveform_sig_rx =884;
8332: waveform_sig_rx =839;
8333: waveform_sig_rx =659;
8334: waveform_sig_rx =800;
8335: waveform_sig_rx =937;
8336: waveform_sig_rx =618;
8337: waveform_sig_rx =718;
8338: waveform_sig_rx =980;
8339: waveform_sig_rx =582;
8340: waveform_sig_rx =773;
8341: waveform_sig_rx =789;
8342: waveform_sig_rx =653;
8343: waveform_sig_rx =808;
8344: waveform_sig_rx =678;
8345: waveform_sig_rx =717;
8346: waveform_sig_rx =595;
8347: waveform_sig_rx =913;
8348: waveform_sig_rx =511;
8349: waveform_sig_rx =713;
8350: waveform_sig_rx =809;
8351: waveform_sig_rx =497;
8352: waveform_sig_rx =699;
8353: waveform_sig_rx =815;
8354: waveform_sig_rx =528;
8355: waveform_sig_rx =586;
8356: waveform_sig_rx =843;
8357: waveform_sig_rx =525;
8358: waveform_sig_rx =548;
8359: waveform_sig_rx =795;
8360: waveform_sig_rx =608;
8361: waveform_sig_rx =422;
8362: waveform_sig_rx =811;
8363: waveform_sig_rx =627;
8364: waveform_sig_rx =474;
8365: waveform_sig_rx =616;
8366: waveform_sig_rx =726;
8367: waveform_sig_rx =466;
8368: waveform_sig_rx =544;
8369: waveform_sig_rx =726;
8370: waveform_sig_rx =498;
8371: waveform_sig_rx =473;
8372: waveform_sig_rx =636;
8373: waveform_sig_rx =636;
8374: waveform_sig_rx =340;
8375: waveform_sig_rx =588;
8376: waveform_sig_rx =713;
8377: waveform_sig_rx =293;
8378: waveform_sig_rx =555;
8379: waveform_sig_rx =699;
8380: waveform_sig_rx =291;
8381: waveform_sig_rx =611;
8382: waveform_sig_rx =435;
8383: waveform_sig_rx =458;
8384: waveform_sig_rx =576;
8385: waveform_sig_rx =400;
8386: waveform_sig_rx =539;
8387: waveform_sig_rx =322;
8388: waveform_sig_rx =636;
8389: waveform_sig_rx =278;
8390: waveform_sig_rx =411;
8391: waveform_sig_rx =594;
8392: waveform_sig_rx =241;
8393: waveform_sig_rx =410;
8394: waveform_sig_rx =573;
8395: waveform_sig_rx =237;
8396: waveform_sig_rx =342;
8397: waveform_sig_rx =577;
8398: waveform_sig_rx =230;
8399: waveform_sig_rx =284;
8400: waveform_sig_rx =549;
8401: waveform_sig_rx =287;
8402: waveform_sig_rx =156;
8403: waveform_sig_rx =539;
8404: waveform_sig_rx =290;
8405: waveform_sig_rx =265;
8406: waveform_sig_rx =336;
8407: waveform_sig_rx =401;
8408: waveform_sig_rx =214;
8409: waveform_sig_rx =209;
8410: waveform_sig_rx =454;
8411: waveform_sig_rx =235;
8412: waveform_sig_rx =124;
8413: waveform_sig_rx =411;
8414: waveform_sig_rx =311;
8415: waveform_sig_rx =49;
8416: waveform_sig_rx =365;
8417: waveform_sig_rx =321;
8418: waveform_sig_rx =28;
8419: waveform_sig_rx =295;
8420: waveform_sig_rx =343;
8421: waveform_sig_rx =60;
8422: waveform_sig_rx =290;
8423: waveform_sig_rx =113;
8424: waveform_sig_rx =240;
8425: waveform_sig_rx =192;
8426: waveform_sig_rx =136;
8427: waveform_sig_rx =238;
8428: waveform_sig_rx =-21;
8429: waveform_sig_rx =387;
8430: waveform_sig_rx =-37;
8431: waveform_sig_rx =132;
8432: waveform_sig_rx =312;
8433: waveform_sig_rx =-105;
8434: waveform_sig_rx =141;
8435: waveform_sig_rx =296;
8436: waveform_sig_rx =-93;
8437: waveform_sig_rx =59;
8438: waveform_sig_rx =310;
8439: waveform_sig_rx =-119;
8440: waveform_sig_rx =42;
8441: waveform_sig_rx =252;
8442: waveform_sig_rx =-45;
8443: waveform_sig_rx =-62;
8444: waveform_sig_rx =206;
8445: waveform_sig_rx =-36;
8446: waveform_sig_rx =-8;
8447: waveform_sig_rx =-35;
8448: waveform_sig_rx =186;
8449: waveform_sig_rx =-90;
8450: waveform_sig_rx =-111;
8451: waveform_sig_rx =243;
8452: waveform_sig_rx =-157;
8453: waveform_sig_rx =-128;
8454: waveform_sig_rx =153;
8455: waveform_sig_rx =-78;
8456: waveform_sig_rx =-171;
8457: waveform_sig_rx =45;
8458: waveform_sig_rx =-8;
8459: waveform_sig_rx =-193;
8460: waveform_sig_rx =-62;
8461: waveform_sig_rx =64;
8462: waveform_sig_rx =-240;
8463: waveform_sig_rx =-72;
8464: waveform_sig_rx =-171;
8465: waveform_sig_rx =-99;
8466: waveform_sig_rx =-133;
8467: waveform_sig_rx =-139;
8468: waveform_sig_rx =-131;
8469: waveform_sig_rx =-297;
8470: waveform_sig_rx =75;
8471: waveform_sig_rx =-400;
8472: waveform_sig_rx =-167;
8473: waveform_sig_rx =13;
8474: waveform_sig_rx =-434;
8475: waveform_sig_rx =-126;
8476: waveform_sig_rx =9;
8477: waveform_sig_rx =-476;
8478: waveform_sig_rx =-163;
8479: waveform_sig_rx =-30;
8480: waveform_sig_rx =-471;
8481: waveform_sig_rx =-194;
8482: waveform_sig_rx =-153;
8483: waveform_sig_rx =-313;
8484: waveform_sig_rx =-373;
8485: waveform_sig_rx =-173;
8486: waveform_sig_rx =-237;
8487: waveform_sig_rx =-403;
8488: waveform_sig_rx =-307;
8489: waveform_sig_rx =-94;
8490: waveform_sig_rx =-501;
8491: waveform_sig_rx =-316;
8492: waveform_sig_rx =-132;
8493: waveform_sig_rx =-472;
8494: waveform_sig_rx =-376;
8495: waveform_sig_rx =-206;
8496: waveform_sig_rx =-372;
8497: waveform_sig_rx =-506;
8498: waveform_sig_rx =-264;
8499: waveform_sig_rx =-292;
8500: waveform_sig_rx =-513;
8501: waveform_sig_rx =-377;
8502: waveform_sig_rx =-235;
8503: waveform_sig_rx =-535;
8504: waveform_sig_rx =-398;
8505: waveform_sig_rx =-407;
8506: waveform_sig_rx =-403;
8507: waveform_sig_rx =-435;
8508: waveform_sig_rx =-380;
8509: waveform_sig_rx =-470;
8510: waveform_sig_rx =-543;
8511: waveform_sig_rx =-216;
8512: waveform_sig_rx =-726;
8513: waveform_sig_rx =-392;
8514: waveform_sig_rx =-333;
8515: waveform_sig_rx =-749;
8516: waveform_sig_rx =-361;
8517: waveform_sig_rx =-381;
8518: waveform_sig_rx =-729;
8519: waveform_sig_rx =-447;
8520: waveform_sig_rx =-377;
8521: waveform_sig_rx =-687;
8522: waveform_sig_rx =-523;
8523: waveform_sig_rx =-441;
8524: waveform_sig_rx =-589;
8525: waveform_sig_rx =-717;
8526: waveform_sig_rx =-414;
8527: waveform_sig_rx =-547;
8528: waveform_sig_rx =-740;
8529: waveform_sig_rx =-560;
8530: waveform_sig_rx =-432;
8531: waveform_sig_rx =-781;
8532: waveform_sig_rx =-565;
8533: waveform_sig_rx =-446;
8534: waveform_sig_rx =-755;
8535: waveform_sig_rx =-668;
8536: waveform_sig_rx =-506;
8537: waveform_sig_rx =-648;
8538: waveform_sig_rx =-773;
8539: waveform_sig_rx =-559;
8540: waveform_sig_rx =-578;
8541: waveform_sig_rx =-801;
8542: waveform_sig_rx =-657;
8543: waveform_sig_rx =-478;
8544: waveform_sig_rx =-854;
8545: waveform_sig_rx =-640;
8546: waveform_sig_rx =-680;
8547: waveform_sig_rx =-724;
8548: waveform_sig_rx =-662;
8549: waveform_sig_rx =-672;
8550: waveform_sig_rx =-782;
8551: waveform_sig_rx =-755;
8552: waveform_sig_rx =-543;
8553: waveform_sig_rx =-968;
8554: waveform_sig_rx =-636;
8555: waveform_sig_rx =-647;
8556: waveform_sig_rx =-929;
8557: waveform_sig_rx =-660;
8558: waveform_sig_rx =-628;
8559: waveform_sig_rx =-945;
8560: waveform_sig_rx =-725;
8561: waveform_sig_rx =-613;
8562: waveform_sig_rx =-956;
8563: waveform_sig_rx =-771;
8564: waveform_sig_rx =-674;
8565: waveform_sig_rx =-837;
8566: waveform_sig_rx =-973;
8567: waveform_sig_rx =-643;
8568: waveform_sig_rx =-822;
8569: waveform_sig_rx =-986;
8570: waveform_sig_rx =-744;
8571: waveform_sig_rx =-711;
8572: waveform_sig_rx =-1008;
8573: waveform_sig_rx =-779;
8574: waveform_sig_rx =-754;
8575: waveform_sig_rx =-926;
8576: waveform_sig_rx =-908;
8577: waveform_sig_rx =-738;
8578: waveform_sig_rx =-829;
8579: waveform_sig_rx =-1074;
8580: waveform_sig_rx =-744;
8581: waveform_sig_rx =-791;
8582: waveform_sig_rx =-1082;
8583: waveform_sig_rx =-819;
8584: waveform_sig_rx =-756;
8585: waveform_sig_rx =-1115;
8586: waveform_sig_rx =-793;
8587: waveform_sig_rx =-971;
8588: waveform_sig_rx =-918;
8589: waveform_sig_rx =-897;
8590: waveform_sig_rx =-926;
8591: waveform_sig_rx =-967;
8592: waveform_sig_rx =-974;
8593: waveform_sig_rx =-785;
8594: waveform_sig_rx =-1146;
8595: waveform_sig_rx =-871;
8596: waveform_sig_rx =-860;
8597: waveform_sig_rx =-1161;
8598: waveform_sig_rx =-889;
8599: waveform_sig_rx =-842;
8600: waveform_sig_rx =-1186;
8601: waveform_sig_rx =-936;
8602: waveform_sig_rx =-826;
8603: waveform_sig_rx =-1161;
8604: waveform_sig_rx =-1005;
8605: waveform_sig_rx =-850;
8606: waveform_sig_rx =-1089;
8607: waveform_sig_rx =-1167;
8608: waveform_sig_rx =-778;
8609: waveform_sig_rx =-1090;
8610: waveform_sig_rx =-1112;
8611: waveform_sig_rx =-961;
8612: waveform_sig_rx =-957;
8613: waveform_sig_rx =-1137;
8614: waveform_sig_rx =-1035;
8615: waveform_sig_rx =-901;
8616: waveform_sig_rx =-1119;
8617: waveform_sig_rx =-1151;
8618: waveform_sig_rx =-843;
8619: waveform_sig_rx =-1089;
8620: waveform_sig_rx =-1243;
8621: waveform_sig_rx =-876;
8622: waveform_sig_rx =-1038;
8623: waveform_sig_rx =-1225;
8624: waveform_sig_rx =-983;
8625: waveform_sig_rx =-953;
8626: waveform_sig_rx =-1249;
8627: waveform_sig_rx =-985;
8628: waveform_sig_rx =-1148;
8629: waveform_sig_rx =-1045;
8630: waveform_sig_rx =-1081;
8631: waveform_sig_rx =-1080;
8632: waveform_sig_rx =-1122;
8633: waveform_sig_rx =-1132;
8634: waveform_sig_rx =-954;
8635: waveform_sig_rx =-1269;
8636: waveform_sig_rx =-1035;
8637: waveform_sig_rx =-998;
8638: waveform_sig_rx =-1281;
8639: waveform_sig_rx =-1047;
8640: waveform_sig_rx =-927;
8641: waveform_sig_rx =-1376;
8642: waveform_sig_rx =-1033;
8643: waveform_sig_rx =-920;
8644: waveform_sig_rx =-1378;
8645: waveform_sig_rx =-1031;
8646: waveform_sig_rx =-1002;
8647: waveform_sig_rx =-1233;
8648: waveform_sig_rx =-1210;
8649: waveform_sig_rx =-970;
8650: waveform_sig_rx =-1195;
8651: waveform_sig_rx =-1206;
8652: waveform_sig_rx =-1106;
8653: waveform_sig_rx =-1026;
8654: waveform_sig_rx =-1289;
8655: waveform_sig_rx =-1144;
8656: waveform_sig_rx =-995;
8657: waveform_sig_rx =-1267;
8658: waveform_sig_rx =-1213;
8659: waveform_sig_rx =-944;
8660: waveform_sig_rx =-1209;
8661: waveform_sig_rx =-1294;
8662: waveform_sig_rx =-962;
8663: waveform_sig_rx =-1149;
8664: waveform_sig_rx =-1282;
8665: waveform_sig_rx =-1060;
8666: waveform_sig_rx =-1057;
8667: waveform_sig_rx =-1303;
8668: waveform_sig_rx =-1065;
8669: waveform_sig_rx =-1248;
8670: waveform_sig_rx =-1068;
8671: waveform_sig_rx =-1198;
8672: waveform_sig_rx =-1124;
8673: waveform_sig_rx =-1174;
8674: waveform_sig_rx =-1228;
8675: waveform_sig_rx =-990;
8676: waveform_sig_rx =-1391;
8677: waveform_sig_rx =-1117;
8678: waveform_sig_rx =-1013;
8679: waveform_sig_rx =-1434;
8680: waveform_sig_rx =-1033;
8681: waveform_sig_rx =-1014;
8682: waveform_sig_rx =-1458;
8683: waveform_sig_rx =-995;
8684: waveform_sig_rx =-1071;
8685: waveform_sig_rx =-1369;
8686: waveform_sig_rx =-1057;
8687: waveform_sig_rx =-1106;
8688: waveform_sig_rx =-1219;
8689: waveform_sig_rx =-1264;
8690: waveform_sig_rx =-997;
8691: waveform_sig_rx =-1186;
8692: waveform_sig_rx =-1273;
8693: waveform_sig_rx =-1105;
8694: waveform_sig_rx =-1049;
8695: waveform_sig_rx =-1325;
8696: waveform_sig_rx =-1127;
8697: waveform_sig_rx =-1026;
8698: waveform_sig_rx =-1286;
8699: waveform_sig_rx =-1226;
8700: waveform_sig_rx =-946;
8701: waveform_sig_rx =-1262;
8702: waveform_sig_rx =-1268;
8703: waveform_sig_rx =-982;
8704: waveform_sig_rx =-1205;
8705: waveform_sig_rx =-1244;
8706: waveform_sig_rx =-1103;
8707: waveform_sig_rx =-1048;
8708: waveform_sig_rx =-1274;
8709: waveform_sig_rx =-1115;
8710: waveform_sig_rx =-1186;
8711: waveform_sig_rx =-1097;
8712: waveform_sig_rx =-1210;
8713: waveform_sig_rx =-1050;
8714: waveform_sig_rx =-1258;
8715: waveform_sig_rx =-1146;
8716: waveform_sig_rx =-950;
8717: waveform_sig_rx =-1411;
8718: waveform_sig_rx =-974;
8719: waveform_sig_rx =-1063;
8720: waveform_sig_rx =-1373;
8721: waveform_sig_rx =-944;
8722: waveform_sig_rx =-1071;
8723: waveform_sig_rx =-1349;
8724: waveform_sig_rx =-987;
8725: waveform_sig_rx =-1054;
8726: waveform_sig_rx =-1289;
8727: waveform_sig_rx =-1043;
8728: waveform_sig_rx =-1017;
8729: waveform_sig_rx =-1195;
8730: waveform_sig_rx =-1206;
8731: waveform_sig_rx =-933;
8732: waveform_sig_rx =-1165;
8733: waveform_sig_rx =-1209;
8734: waveform_sig_rx =-1045;
8735: waveform_sig_rx =-973;
8736: waveform_sig_rx =-1304;
8737: waveform_sig_rx =-1028;
8738: waveform_sig_rx =-965;
8739: waveform_sig_rx =-1264;
8740: waveform_sig_rx =-1070;
8741: waveform_sig_rx =-954;
8742: waveform_sig_rx =-1163;
8743: waveform_sig_rx =-1152;
8744: waveform_sig_rx =-966;
8745: waveform_sig_rx =-1056;
8746: waveform_sig_rx =-1214;
8747: waveform_sig_rx =-1020;
8748: waveform_sig_rx =-931;
8749: waveform_sig_rx =-1257;
8750: waveform_sig_rx =-949;
8751: waveform_sig_rx =-1113;
8752: waveform_sig_rx =-1026;
8753: waveform_sig_rx =-1069;
8754: waveform_sig_rx =-977;
8755: waveform_sig_rx =-1176;
8756: waveform_sig_rx =-994;
8757: waveform_sig_rx =-925;
8758: waveform_sig_rx =-1279;
8759: waveform_sig_rx =-855;
8760: waveform_sig_rx =-1023;
8761: waveform_sig_rx =-1216;
8762: waveform_sig_rx =-856;
8763: waveform_sig_rx =-985;
8764: waveform_sig_rx =-1200;
8765: waveform_sig_rx =-878;
8766: waveform_sig_rx =-932;
8767: waveform_sig_rx =-1160;
8768: waveform_sig_rx =-937;
8769: waveform_sig_rx =-878;
8770: waveform_sig_rx =-1084;
8771: waveform_sig_rx =-1070;
8772: waveform_sig_rx =-803;
8773: waveform_sig_rx =-1029;
8774: waveform_sig_rx =-1075;
8775: waveform_sig_rx =-875;
8776: waveform_sig_rx =-882;
8777: waveform_sig_rx =-1176;
8778: waveform_sig_rx =-818;
8779: waveform_sig_rx =-890;
8780: waveform_sig_rx =-1067;
8781: waveform_sig_rx =-920;
8782: waveform_sig_rx =-824;
8783: waveform_sig_rx =-950;
8784: waveform_sig_rx =-1074;
8785: waveform_sig_rx =-768;
8786: waveform_sig_rx =-900;
8787: waveform_sig_rx =-1112;
8788: waveform_sig_rx =-766;
8789: waveform_sig_rx =-845;
8790: waveform_sig_rx =-1085;
8791: waveform_sig_rx =-753;
8792: waveform_sig_rx =-1030;
8793: waveform_sig_rx =-812;
8794: waveform_sig_rx =-938;
8795: waveform_sig_rx =-827;
8796: waveform_sig_rx =-1009;
8797: waveform_sig_rx =-833;
8798: waveform_sig_rx =-765;
8799: waveform_sig_rx =-1088;
8800: waveform_sig_rx =-675;
8801: waveform_sig_rx =-866;
8802: waveform_sig_rx =-1010;
8803: waveform_sig_rx =-692;
8804: waveform_sig_rx =-823;
8805: waveform_sig_rx =-995;
8806: waveform_sig_rx =-747;
8807: waveform_sig_rx =-738;
8808: waveform_sig_rx =-999;
8809: waveform_sig_rx =-781;
8810: waveform_sig_rx =-661;
8811: waveform_sig_rx =-973;
8812: waveform_sig_rx =-856;
8813: waveform_sig_rx =-592;
8814: waveform_sig_rx =-908;
8815: waveform_sig_rx =-846;
8816: waveform_sig_rx =-690;
8817: waveform_sig_rx =-710;
8818: waveform_sig_rx =-929;
8819: waveform_sig_rx =-661;
8820: waveform_sig_rx =-684;
8821: waveform_sig_rx =-859;
8822: waveform_sig_rx =-766;
8823: waveform_sig_rx =-591;
8824: waveform_sig_rx =-776;
8825: waveform_sig_rx =-892;
8826: waveform_sig_rx =-523;
8827: waveform_sig_rx =-766;
8828: waveform_sig_rx =-901;
8829: waveform_sig_rx =-527;
8830: waveform_sig_rx =-705;
8831: waveform_sig_rx =-833;
8832: waveform_sig_rx =-571;
8833: waveform_sig_rx =-852;
8834: waveform_sig_rx =-556;
8835: waveform_sig_rx =-748;
8836: waveform_sig_rx =-599;
8837: waveform_sig_rx =-765;
8838: waveform_sig_rx =-632;
8839: waveform_sig_rx =-557;
8840: waveform_sig_rx =-851;
8841: waveform_sig_rx =-479;
8842: waveform_sig_rx =-623;
8843: waveform_sig_rx =-800;
8844: waveform_sig_rx =-456;
8845: waveform_sig_rx =-564;
8846: waveform_sig_rx =-812;
8847: waveform_sig_rx =-477;
8848: waveform_sig_rx =-496;
8849: waveform_sig_rx =-795;
8850: waveform_sig_rx =-489;
8851: waveform_sig_rx =-444;
8852: waveform_sig_rx =-776;
8853: waveform_sig_rx =-553;
8854: waveform_sig_rx =-395;
8855: waveform_sig_rx =-664;
8856: waveform_sig_rx =-582;
8857: waveform_sig_rx =-477;
8858: waveform_sig_rx =-451;
8859: waveform_sig_rx =-694;
8860: waveform_sig_rx =-456;
8861: waveform_sig_rx =-414;
8862: waveform_sig_rx =-649;
8863: waveform_sig_rx =-526;
8864: waveform_sig_rx =-303;
8865: waveform_sig_rx =-599;
8866: waveform_sig_rx =-598;
8867: waveform_sig_rx =-249;
8868: waveform_sig_rx =-557;
8869: waveform_sig_rx =-582;
8870: waveform_sig_rx =-304;
8871: waveform_sig_rx =-440;
8872: waveform_sig_rx =-531;
8873: waveform_sig_rx =-361;
8874: waveform_sig_rx =-548;
8875: waveform_sig_rx =-318;
8876: waveform_sig_rx =-517;
8877: waveform_sig_rx =-293;
8878: waveform_sig_rx =-527;
8879: waveform_sig_rx =-352;
8880: waveform_sig_rx =-271;
8881: waveform_sig_rx =-604;
8882: waveform_sig_rx =-196;
8883: waveform_sig_rx =-357;
8884: waveform_sig_rx =-546;
8885: waveform_sig_rx =-174;
8886: waveform_sig_rx =-306;
8887: waveform_sig_rx =-565;
8888: waveform_sig_rx =-157;
8889: waveform_sig_rx =-250;
8890: waveform_sig_rx =-540;
8891: waveform_sig_rx =-174;
8892: waveform_sig_rx =-237;
8893: waveform_sig_rx =-472;
8894: waveform_sig_rx =-238;
8895: waveform_sig_rx =-190;
8896: waveform_sig_rx =-338;
8897: waveform_sig_rx =-330;
8898: waveform_sig_rx =-213;
8899: waveform_sig_rx =-120;
8900: waveform_sig_rx =-482;
8901: waveform_sig_rx =-120;
8902: waveform_sig_rx =-133;
8903: waveform_sig_rx =-426;
8904: waveform_sig_rx =-150;
8905: waveform_sig_rx =-64;
8906: waveform_sig_rx =-322;
8907: waveform_sig_rx =-246;
8908: waveform_sig_rx =-32;
8909: waveform_sig_rx =-247;
8910: waveform_sig_rx =-289;
8911: waveform_sig_rx =-47;
8912: waveform_sig_rx =-157;
8913: waveform_sig_rx =-269;
8914: waveform_sig_rx =-80;
8915: waveform_sig_rx =-224;
8916: waveform_sig_rx =-23;
8917: waveform_sig_rx =-230;
8918: waveform_sig_rx =24;
8919: waveform_sig_rx =-264;
8920: waveform_sig_rx =-38;
8921: waveform_sig_rx =-9;
8922: waveform_sig_rx =-322;
8923: waveform_sig_rx =107;
8924: waveform_sig_rx =-78;
8925: waveform_sig_rx =-290;
8926: waveform_sig_rx =182;
8927: waveform_sig_rx =-59;
8928: waveform_sig_rx =-271;
8929: waveform_sig_rx =209;
8930: waveform_sig_rx =-51;
8931: waveform_sig_rx =-175;
8932: waveform_sig_rx =122;
8933: waveform_sig_rx =23;
8934: waveform_sig_rx =-102;
8935: waveform_sig_rx =-19;
8936: waveform_sig_rx =125;
8937: waveform_sig_rx =-16;
8938: waveform_sig_rx =-99;
8939: waveform_sig_rx =163;
8940: waveform_sig_rx =98;
8941: waveform_sig_rx =-185;
8942: waveform_sig_rx =235;
8943: waveform_sig_rx =87;
8944: waveform_sig_rx =-74;
8945: waveform_sig_rx =122;
8946: waveform_sig_rx =196;
8947: waveform_sig_rx =4;
8948: waveform_sig_rx =32;
8949: waveform_sig_rx =272;
8950: waveform_sig_rx =42;
8951: waveform_sig_rx =16;
8952: waveform_sig_rx =259;
8953: waveform_sig_rx =150;
8954: waveform_sig_rx =43;
8955: waveform_sig_rx =215;
8956: waveform_sig_rx =87;
8957: waveform_sig_rx =229;
8958: waveform_sig_rx =74;
8959: waveform_sig_rx =313;
8960: waveform_sig_rx =-27;
8961: waveform_sig_rx =317;
8962: waveform_sig_rx =240;
8963: waveform_sig_rx =-52;
8964: waveform_sig_rx =477;
8965: waveform_sig_rx =130;
8966: waveform_sig_rx =61;
8967: waveform_sig_rx =473;
8968: waveform_sig_rx =167;
8969: waveform_sig_rx =104;
8970: waveform_sig_rx =405;
8971: waveform_sig_rx =264;
8972: waveform_sig_rx =130;
8973: waveform_sig_rx =347;
8974: waveform_sig_rx =386;
8975: waveform_sig_rx =121;
8976: waveform_sig_rx =268;
8977: waveform_sig_rx =481;
8978: waveform_sig_rx =201;
8979: waveform_sig_rx =249;
8980: waveform_sig_rx =452;
8981: waveform_sig_rx =349;
8982: waveform_sig_rx =145;
8983: waveform_sig_rx =506;
8984: waveform_sig_rx =379;
8985: waveform_sig_rx =198;
8986: waveform_sig_rx =411;
8987: waveform_sig_rx =465;
8988: waveform_sig_rx =264;
8989: waveform_sig_rx =315;
8990: waveform_sig_rx =535;
8991: waveform_sig_rx =345;
8992: waveform_sig_rx =256;
8993: waveform_sig_rx =566;
8994: waveform_sig_rx =459;
8995: waveform_sig_rx =282;
8996: waveform_sig_rx =551;
8997: waveform_sig_rx =351;
8998: waveform_sig_rx =495;
8999: waveform_sig_rx =418;
9000: waveform_sig_rx =515;
9001: waveform_sig_rx =283;
9002: waveform_sig_rx =642;
9003: waveform_sig_rx =449;
9004: waveform_sig_rx =333;
9005: waveform_sig_rx =710;
9006: waveform_sig_rx =395;
9007: waveform_sig_rx =398;
9008: waveform_sig_rx =677;
9009: waveform_sig_rx =498;
9010: waveform_sig_rx =340;
9011: waveform_sig_rx =712;
9012: waveform_sig_rx =552;
9013: waveform_sig_rx =392;
9014: waveform_sig_rx =648;
9015: waveform_sig_rx =647;
9016: waveform_sig_rx =413;
9017: waveform_sig_rx =566;
9018: waveform_sig_rx =747;
9019: waveform_sig_rx =452;
9020: waveform_sig_rx =519;
9021: waveform_sig_rx =747;
9022: waveform_sig_rx =575;
9023: waveform_sig_rx =449;
9024: waveform_sig_rx =758;
9025: waveform_sig_rx =616;
9026: waveform_sig_rx =504;
9027: waveform_sig_rx =658;
9028: waveform_sig_rx =755;
9029: waveform_sig_rx =538;
9030: waveform_sig_rx =553;
9031: waveform_sig_rx =847;
9032: waveform_sig_rx =564;
9033: waveform_sig_rx =517;
9034: waveform_sig_rx =878;
9035: waveform_sig_rx =636;
9036: waveform_sig_rx =565;
9037: waveform_sig_rx =822;
9038: waveform_sig_rx =546;
9039: waveform_sig_rx =797;
9040: waveform_sig_rx =652;
9041: waveform_sig_rx =753;
9042: waveform_sig_rx =590;
9043: waveform_sig_rx =844;
9044: waveform_sig_rx =718;
9045: waveform_sig_rx =582;
9046: waveform_sig_rx =916;
9047: waveform_sig_rx =707;
9048: waveform_sig_rx =596;
9049: waveform_sig_rx =970;
9050: waveform_sig_rx =727;
9051: waveform_sig_rx =560;
9052: waveform_sig_rx =984;
9053: waveform_sig_rx =740;
9054: waveform_sig_rx =628;
9055: waveform_sig_rx =891;
9056: waveform_sig_rx =858;
9057: waveform_sig_rx =624;
9058: waveform_sig_rx =823;
9059: waveform_sig_rx =970;
9060: waveform_sig_rx =640;
9061: waveform_sig_rx =801;
9062: waveform_sig_rx =922;
9063: waveform_sig_rx =797;
9064: waveform_sig_rx =737;
9065: waveform_sig_rx =904;
9066: waveform_sig_rx =904;
9067: waveform_sig_rx =703;
9068: waveform_sig_rx =867;
9069: waveform_sig_rx =1071;
9070: waveform_sig_rx =653;
9071: waveform_sig_rx =869;
9072: waveform_sig_rx =1075;
9073: waveform_sig_rx =721;
9074: waveform_sig_rx =819;
9075: waveform_sig_rx =1023;
9076: waveform_sig_rx =865;
9077: waveform_sig_rx =818;
9078: waveform_sig_rx =974;
9079: waveform_sig_rx =806;
9080: waveform_sig_rx =1014;
9081: waveform_sig_rx =837;
9082: waveform_sig_rx =993;
9083: waveform_sig_rx =782;
9084: waveform_sig_rx =1063;
9085: waveform_sig_rx =912;
9086: waveform_sig_rx =782;
9087: waveform_sig_rx =1113;
9088: waveform_sig_rx =884;
9089: waveform_sig_rx =778;
9090: waveform_sig_rx =1156;
9091: waveform_sig_rx =914;
9092: waveform_sig_rx =730;
9093: waveform_sig_rx =1227;
9094: waveform_sig_rx =890;
9095: waveform_sig_rx =818;
9096: waveform_sig_rx =1143;
9097: waveform_sig_rx =990;
9098: waveform_sig_rx =818;
9099: waveform_sig_rx =1069;
9100: waveform_sig_rx =1077;
9101: waveform_sig_rx =881;
9102: waveform_sig_rx =973;
9103: waveform_sig_rx =1112;
9104: waveform_sig_rx =1025;
9105: waveform_sig_rx =852;
9106: waveform_sig_rx =1134;
9107: waveform_sig_rx =1081;
9108: waveform_sig_rx =826;
9109: waveform_sig_rx =1106;
9110: waveform_sig_rx =1167;
9111: waveform_sig_rx =827;
9112: waveform_sig_rx =1062;
9113: waveform_sig_rx =1168;
9114: waveform_sig_rx =908;
9115: waveform_sig_rx =983;
9116: waveform_sig_rx =1163;
9117: waveform_sig_rx =1004;
9118: waveform_sig_rx =989;
9119: waveform_sig_rx =1110;
9120: waveform_sig_rx =972;
9121: waveform_sig_rx =1154;
9122: waveform_sig_rx =976;
9123: waveform_sig_rx =1173;
9124: waveform_sig_rx =892;
9125: waveform_sig_rx =1232;
9126: waveform_sig_rx =1070;
9127: waveform_sig_rx =904;
9128: waveform_sig_rx =1309;
9129: waveform_sig_rx =982;
9130: waveform_sig_rx =920;
9131: waveform_sig_rx =1382;
9132: waveform_sig_rx =957;
9133: waveform_sig_rx =910;
9134: waveform_sig_rx =1368;
9135: waveform_sig_rx =957;
9136: waveform_sig_rx =1025;
9137: waveform_sig_rx =1229;
9138: waveform_sig_rx =1107;
9139: waveform_sig_rx =989;
9140: waveform_sig_rx =1148;
9141: waveform_sig_rx =1211;
9142: waveform_sig_rx =1019;
9143: waveform_sig_rx =1055;
9144: waveform_sig_rx =1263;
9145: waveform_sig_rx =1099;
9146: waveform_sig_rx =969;
9147: waveform_sig_rx =1280;
9148: waveform_sig_rx =1120;
9149: waveform_sig_rx =947;
9150: waveform_sig_rx =1228;
9151: waveform_sig_rx =1202;
9152: waveform_sig_rx =953;
9153: waveform_sig_rx =1173;
9154: waveform_sig_rx =1236;
9155: waveform_sig_rx =1038;
9156: waveform_sig_rx =1074;
9157: waveform_sig_rx =1269;
9158: waveform_sig_rx =1103;
9159: waveform_sig_rx =1044;
9160: waveform_sig_rx =1198;
9161: waveform_sig_rx =1080;
9162: waveform_sig_rx =1181;
9163: waveform_sig_rx =1077;
9164: waveform_sig_rx =1245;
9165: waveform_sig_rx =917;
9166: waveform_sig_rx =1348;
9167: waveform_sig_rx =1053;
9168: waveform_sig_rx =972;
9169: waveform_sig_rx =1407;
9170: waveform_sig_rx =961;
9171: waveform_sig_rx =1056;
9172: waveform_sig_rx =1391;
9173: waveform_sig_rx =974;
9174: waveform_sig_rx =1042;
9175: waveform_sig_rx =1369;
9176: waveform_sig_rx =1029;
9177: waveform_sig_rx =1086;
9178: waveform_sig_rx =1258;
9179: waveform_sig_rx =1187;
9180: waveform_sig_rx =998;
9181: waveform_sig_rx =1215;
9182: waveform_sig_rx =1265;
9183: waveform_sig_rx =1026;
9184: waveform_sig_rx =1077;
9185: waveform_sig_rx =1325;
9186: waveform_sig_rx =1088;
9187: waveform_sig_rx =989;
9188: waveform_sig_rx =1358;
9189: waveform_sig_rx =1100;
9190: waveform_sig_rx =1018;
9191: waveform_sig_rx =1264;
9192: waveform_sig_rx =1200;
9193: waveform_sig_rx =1029;
9194: waveform_sig_rx =1168;
9195: waveform_sig_rx =1267;
9196: waveform_sig_rx =1068;
9197: waveform_sig_rx =1036;
9198: waveform_sig_rx =1348;
9199: waveform_sig_rx =1086;
9200: waveform_sig_rx =1047;
9201: waveform_sig_rx =1250;
9202: waveform_sig_rx =1030;
9203: waveform_sig_rx =1216;
9204: waveform_sig_rx =1120;
9205: waveform_sig_rx =1190;
9206: waveform_sig_rx =982;
9207: waveform_sig_rx =1355;
9208: waveform_sig_rx =1001;
9209: waveform_sig_rx =1036;
9210: waveform_sig_rx =1328;
9211: waveform_sig_rx =934;
9212: waveform_sig_rx =1086;
9213: waveform_sig_rx =1327;
9214: waveform_sig_rx =964;
9215: waveform_sig_rx =1045;
9216: waveform_sig_rx =1320;
9217: waveform_sig_rx =1035;
9218: waveform_sig_rx =1068;
9219: waveform_sig_rx =1206;
9220: waveform_sig_rx =1186;
9221: waveform_sig_rx =906;
9222: waveform_sig_rx =1161;
9223: waveform_sig_rx =1231;
9224: waveform_sig_rx =935;
9225: waveform_sig_rx =1103;
9226: waveform_sig_rx =1278;
9227: waveform_sig_rx =992;
9228: waveform_sig_rx =1021;
9229: waveform_sig_rx =1255;
9230: waveform_sig_rx =1050;
9231: waveform_sig_rx =1002;
9232: waveform_sig_rx =1169;
9233: waveform_sig_rx =1200;
9234: waveform_sig_rx =951;
9235: waveform_sig_rx =1081;
9236: waveform_sig_rx =1249;
9237: waveform_sig_rx =949;
9238: waveform_sig_rx =1002;
9239: waveform_sig_rx =1292;
9240: waveform_sig_rx =977;
9241: waveform_sig_rx =1044;
9242: waveform_sig_rx =1162;
9243: waveform_sig_rx =962;
9244: waveform_sig_rx =1181;
9245: waveform_sig_rx =1028;
9246: waveform_sig_rx =1107;
9247: waveform_sig_rx =928;
9248: waveform_sig_rx =1266;
9249: waveform_sig_rx =908;
9250: waveform_sig_rx =998;
9251: waveform_sig_rx =1224;
9252: waveform_sig_rx =870;
9253: waveform_sig_rx =1018;
9254: waveform_sig_rx =1221;
9255: waveform_sig_rx =920;
9256: waveform_sig_rx =951;
9257: waveform_sig_rx =1217;
9258: waveform_sig_rx =954;
9259: waveform_sig_rx =917;
9260: waveform_sig_rx =1152;
9261: waveform_sig_rx =1062;
9262: waveform_sig_rx =790;
9263: waveform_sig_rx =1160;
9264: waveform_sig_rx =1057;
9265: waveform_sig_rx =865;
9266: waveform_sig_rx =1015;
9267: waveform_sig_rx =1119;
9268: waveform_sig_rx =919;
9269: waveform_sig_rx =932;
9270: waveform_sig_rx =1129;
9271: waveform_sig_rx =964;
9272: waveform_sig_rx =878;
9273: waveform_sig_rx =1047;
9274: waveform_sig_rx =1093;
9275: waveform_sig_rx =786;
9276: waveform_sig_rx =979;
9277: waveform_sig_rx =1142;
9278: waveform_sig_rx =758;
9279: waveform_sig_rx =928;
9280: waveform_sig_rx =1132;
9281: waveform_sig_rx =792;
9282: waveform_sig_rx =959;
9283: waveform_sig_rx =943;
9284: waveform_sig_rx =857;
9285: waveform_sig_rx =1033;
9286: waveform_sig_rx =839;
9287: waveform_sig_rx =1012;
9288: waveform_sig_rx =767;
9289: waveform_sig_rx =1116;
9290: waveform_sig_rx =787;
9291: waveform_sig_rx =836;
9292: waveform_sig_rx =1086;
9293: waveform_sig_rx =747;
9294: waveform_sig_rx =851;
9295: waveform_sig_rx =1095;
9296: waveform_sig_rx =764;
9297: waveform_sig_rx =755;
9298: waveform_sig_rx =1094;
9299: waveform_sig_rx =753;
9300: waveform_sig_rx =751;
9301: waveform_sig_rx =1041;
9302: waveform_sig_rx =839;
9303: waveform_sig_rx =646;
9304: waveform_sig_rx =1000;
9305: waveform_sig_rx =849;
9306: waveform_sig_rx =736;
9307: waveform_sig_rx =817;
9308: waveform_sig_rx =934;
9309: waveform_sig_rx =764;
9310: waveform_sig_rx =705;
9311: waveform_sig_rx =974;
9312: waveform_sig_rx =760;
9313: waveform_sig_rx =659;
9314: waveform_sig_rx =918;
9315: waveform_sig_rx =864;
9316: waveform_sig_rx =591;
9317: waveform_sig_rx =851;
9318: waveform_sig_rx =921;
9319: waveform_sig_rx =571;
9320: waveform_sig_rx =791;
9321: waveform_sig_rx =898;
9322: waveform_sig_rx =626;
9323: waveform_sig_rx =784;
9324: waveform_sig_rx =702;
9325: waveform_sig_rx =731;
9326: waveform_sig_rx =792;
9327: waveform_sig_rx =642;
9328: waveform_sig_rx =830;
9329: waveform_sig_rx =515;
9330: waveform_sig_rx =927;
9331: waveform_sig_rx =572;
9332: waveform_sig_rx =613;
9333: waveform_sig_rx =891;
9334: waveform_sig_rx =507;
9335: waveform_sig_rx =654;
9336: waveform_sig_rx =898;
9337: waveform_sig_rx =518;
9338: waveform_sig_rx =565;
9339: waveform_sig_rx =898;
9340: waveform_sig_rx =515;
9341: waveform_sig_rx =537;
9342: waveform_sig_rx =833;
9343: waveform_sig_rx =545;
9344: waveform_sig_rx =471;
9345: waveform_sig_rx =763;
9346: waveform_sig_rx =579;
9347: waveform_sig_rx =568;
9348: waveform_sig_rx =519;
9349: waveform_sig_rx =735;
9350: waveform_sig_rx =518;
9351: waveform_sig_rx =428;
9352: waveform_sig_rx =827;
9353: waveform_sig_rx =458;
9354: waveform_sig_rx =447;
9355: waveform_sig_rx =715;
9356: waveform_sig_rx =558;
9357: waveform_sig_rx =385;
9358: waveform_sig_rx =592;
9359: waveform_sig_rx =638;
9360: waveform_sig_rx =361;
9361: waveform_sig_rx =496;
9362: waveform_sig_rx =675;
9363: waveform_sig_rx =388;
9364: waveform_sig_rx =521;
9365: waveform_sig_rx =461;
9366: waveform_sig_rx =467;
9367: waveform_sig_rx =489;
9368: waveform_sig_rx =423;
9369: waveform_sig_rx =542;
9370: waveform_sig_rx =258;
9371: waveform_sig_rx =682;
9372: waveform_sig_rx =278;
9373: waveform_sig_rx =372;
9374: waveform_sig_rx =651;
9375: waveform_sig_rx =192;
9376: waveform_sig_rx =411;
9377: waveform_sig_rx =635;
9378: waveform_sig_rx =185;
9379: waveform_sig_rx =367;
9380: waveform_sig_rx =582;
9381: waveform_sig_rx =176;
9382: waveform_sig_rx =351;
9383: waveform_sig_rx =479;
9384: waveform_sig_rx =334;
9385: waveform_sig_rx =225;
9386: waveform_sig_rx =435;
9387: waveform_sig_rx =388;
9388: waveform_sig_rx =216;
9389: waveform_sig_rx =264;
9390: waveform_sig_rx =514;
9391: waveform_sig_rx =144;
9392: waveform_sig_rx =219;
9393: waveform_sig_rx =493;
9394: waveform_sig_rx =145;
9395: waveform_sig_rx =215;
9396: waveform_sig_rx =377;
9397: waveform_sig_rx =281;
9398: waveform_sig_rx =100;
9399: waveform_sig_rx =302;
9400: waveform_sig_rx =345;
9401: waveform_sig_rx =68;
9402: waveform_sig_rx =199;
9403: waveform_sig_rx =367;
9404: waveform_sig_rx =96;
9405: waveform_sig_rx =207;
9406: waveform_sig_rx =171;
9407: waveform_sig_rx =190;
9408: waveform_sig_rx =178;
9409: waveform_sig_rx =173;
9410: waveform_sig_rx =191;
9411: waveform_sig_rx =-11;
9412: waveform_sig_rx =417;
9413: waveform_sig_rx =-89;
9414: waveform_sig_rx =130;
9415: waveform_sig_rx =342;
9416: waveform_sig_rx =-130;
9417: waveform_sig_rx =194;
9418: waveform_sig_rx =267;
9419: waveform_sig_rx =-96;
9420: waveform_sig_rx =130;
9421: waveform_sig_rx =216;
9422: waveform_sig_rx =-34;
9423: waveform_sig_rx =42;
9424: waveform_sig_rx =171;
9425: waveform_sig_rx =77;
9426: waveform_sig_rx =-156;
9427: waveform_sig_rx =204;
9428: waveform_sig_rx =80;
9429: waveform_sig_rx =-127;
9430: waveform_sig_rx =33;
9431: waveform_sig_rx =157;
9432: waveform_sig_rx =-148;
9433: waveform_sig_rx =-21;
9434: waveform_sig_rx =160;
9435: waveform_sig_rx =-93;
9436: waveform_sig_rx =-116;
9437: waveform_sig_rx =95;
9438: waveform_sig_rx =-17;
9439: waveform_sig_rx =-214;
9440: waveform_sig_rx =22;
9441: waveform_sig_rx =35;
9442: waveform_sig_rx =-197;
9443: waveform_sig_rx =-112;
9444: waveform_sig_rx =100;
9445: waveform_sig_rx =-242;
9446: waveform_sig_rx =-91;
9447: waveform_sig_rx =-61;
9448: waveform_sig_rx =-169;
9449: waveform_sig_rx =-75;
9450: waveform_sig_rx =-88;
9451: waveform_sig_rx =-186;
9452: waveform_sig_rx =-214;
9453: waveform_sig_rx =51;
9454: waveform_sig_rx =-410;
9455: waveform_sig_rx =-94;
9456: waveform_sig_rx =-85;
9457: waveform_sig_rx =-364;
9458: waveform_sig_rx =-156;
9459: waveform_sig_rx =-75;
9460: waveform_sig_rx =-350;
9461: waveform_sig_rx =-278;
9462: waveform_sig_rx =-19;
9463: waveform_sig_rx =-395;
9464: waveform_sig_rx =-281;
9465: waveform_sig_rx =-110;
9466: waveform_sig_rx =-302;
9467: waveform_sig_rx =-426;
9468: waveform_sig_rx =-93;
9469: waveform_sig_rx =-257;
9470: waveform_sig_rx =-400;
9471: waveform_sig_rx =-248;
9472: waveform_sig_rx =-156;
9473: waveform_sig_rx =-446;
9474: waveform_sig_rx =-298;
9475: waveform_sig_rx =-180;
9476: waveform_sig_rx =-424;
9477: waveform_sig_rx =-393;
9478: waveform_sig_rx =-249;
9479: waveform_sig_rx =-273;
9480: waveform_sig_rx =-541;
9481: waveform_sig_rx =-291;
9482: waveform_sig_rx =-215;
9483: waveform_sig_rx =-593;
9484: waveform_sig_rx =-344;
9485: waveform_sig_rx =-205;
9486: waveform_sig_rx =-596;
9487: waveform_sig_rx =-305;
9488: waveform_sig_rx =-442;
9489: waveform_sig_rx =-451;
9490: waveform_sig_rx =-352;
9491: waveform_sig_rx =-462;
9492: waveform_sig_rx =-429;
9493: waveform_sig_rx =-528;
9494: waveform_sig_rx =-279;
9495: waveform_sig_rx =-619;
9496: waveform_sig_rx =-446;
9497: waveform_sig_rx =-360;
9498: waveform_sig_rx =-633;
9499: waveform_sig_rx =-467;
9500: waveform_sig_rx =-297;
9501: waveform_sig_rx =-693;
9502: waveform_sig_rx =-535;
9503: waveform_sig_rx =-287;
9504: waveform_sig_rx =-704;
9505: waveform_sig_rx =-542;
9506: waveform_sig_rx =-388;
9507: waveform_sig_rx =-569;
9508: waveform_sig_rx =-701;
9509: waveform_sig_rx =-354;
9510: waveform_sig_rx =-569;
9511: waveform_sig_rx =-709;
9512: waveform_sig_rx =-513;
9513: waveform_sig_rx =-480;
9514: waveform_sig_rx =-698;
9515: waveform_sig_rx =-610;
9516: waveform_sig_rx =-495;
9517: waveform_sig_rx =-619;
9518: waveform_sig_rx =-756;
9519: waveform_sig_rx =-471;
9520: waveform_sig_rx =-567;
9521: waveform_sig_rx =-869;
9522: waveform_sig_rx =-488;
9523: waveform_sig_rx =-594;
9524: waveform_sig_rx =-854;
9525: waveform_sig_rx =-599;
9526: waveform_sig_rx =-570;
9527: waveform_sig_rx =-824;
9528: waveform_sig_rx =-609;
9529: waveform_sig_rx =-775;
9530: waveform_sig_rx =-656;
9531: waveform_sig_rx =-694;
9532: waveform_sig_rx =-709;
9533: waveform_sig_rx =-683;
9534: waveform_sig_rx =-822;
9535: waveform_sig_rx =-510;
9536: waveform_sig_rx =-902;
9537: waveform_sig_rx =-706;
9538: waveform_sig_rx =-565;
9539: waveform_sig_rx =-927;
9540: waveform_sig_rx =-715;
9541: waveform_sig_rx =-546;
9542: waveform_sig_rx =-973;
9543: waveform_sig_rx =-766;
9544: waveform_sig_rx =-558;
9545: waveform_sig_rx =-987;
9546: waveform_sig_rx =-789;
9547: waveform_sig_rx =-624;
9548: waveform_sig_rx =-885;
9549: waveform_sig_rx =-951;
9550: waveform_sig_rx =-609;
9551: waveform_sig_rx =-866;
9552: waveform_sig_rx =-893;
9553: waveform_sig_rx =-811;
9554: waveform_sig_rx =-711;
9555: waveform_sig_rx =-933;
9556: waveform_sig_rx =-901;
9557: waveform_sig_rx =-662;
9558: waveform_sig_rx =-935;
9559: waveform_sig_rx =-995;
9560: waveform_sig_rx =-631;
9561: waveform_sig_rx =-909;
9562: waveform_sig_rx =-1038;
9563: waveform_sig_rx =-701;
9564: waveform_sig_rx =-871;
9565: waveform_sig_rx =-1003;
9566: waveform_sig_rx =-859;
9567: waveform_sig_rx =-768;
9568: waveform_sig_rx =-1033;
9569: waveform_sig_rx =-866;
9570: waveform_sig_rx =-955;
9571: waveform_sig_rx =-890;
9572: waveform_sig_rx =-922;
9573: waveform_sig_rx =-887;
9574: waveform_sig_rx =-922;
9575: waveform_sig_rx =-1042;
9576: waveform_sig_rx =-718;
9577: waveform_sig_rx =-1144;
9578: waveform_sig_rx =-926;
9579: waveform_sig_rx =-757;
9580: waveform_sig_rx =-1208;
9581: waveform_sig_rx =-912;
9582: waveform_sig_rx =-759;
9583: waveform_sig_rx =-1249;
9584: waveform_sig_rx =-884;
9585: waveform_sig_rx =-806;
9586: waveform_sig_rx =-1218;
9587: waveform_sig_rx =-913;
9588: waveform_sig_rx =-910;
9589: waveform_sig_rx =-1041;
9590: waveform_sig_rx =-1129;
9591: waveform_sig_rx =-864;
9592: waveform_sig_rx =-1016;
9593: waveform_sig_rx =-1122;
9594: waveform_sig_rx =-984;
9595: waveform_sig_rx =-863;
9596: waveform_sig_rx =-1174;
9597: waveform_sig_rx =-1033;
9598: waveform_sig_rx =-829;
9599: waveform_sig_rx =-1162;
9600: waveform_sig_rx =-1119;
9601: waveform_sig_rx =-820;
9602: waveform_sig_rx =-1116;
9603: waveform_sig_rx =-1173;
9604: waveform_sig_rx =-909;
9605: waveform_sig_rx =-1062;
9606: waveform_sig_rx =-1162;
9607: waveform_sig_rx =-1060;
9608: waveform_sig_rx =-918;
9609: waveform_sig_rx =-1214;
9610: waveform_sig_rx =-1056;
9611: waveform_sig_rx =-1085;
9612: waveform_sig_rx =-1071;
9613: waveform_sig_rx =-1115;
9614: waveform_sig_rx =-1032;
9615: waveform_sig_rx =-1140;
9616: waveform_sig_rx =-1146;
9617: waveform_sig_rx =-876;
9618: waveform_sig_rx =-1332;
9619: waveform_sig_rx =-1010;
9620: waveform_sig_rx =-963;
9621: waveform_sig_rx =-1348;
9622: waveform_sig_rx =-970;
9623: waveform_sig_rx =-950;
9624: waveform_sig_rx =-1367;
9625: waveform_sig_rx =-996;
9626: waveform_sig_rx =-991;
9627: waveform_sig_rx =-1311;
9628: waveform_sig_rx =-1056;
9629: waveform_sig_rx =-1044;
9630: waveform_sig_rx =-1141;
9631: waveform_sig_rx =-1252;
9632: waveform_sig_rx =-958;
9633: waveform_sig_rx =-1125;
9634: waveform_sig_rx =-1272;
9635: waveform_sig_rx =-1062;
9636: waveform_sig_rx =-1002;
9637: waveform_sig_rx =-1316;
9638: waveform_sig_rx =-1100;
9639: waveform_sig_rx =-995;
9640: waveform_sig_rx =-1280;
9641: waveform_sig_rx =-1171;
9642: waveform_sig_rx =-990;
9643: waveform_sig_rx =-1190;
9644: waveform_sig_rx =-1267;
9645: waveform_sig_rx =-1035;
9646: waveform_sig_rx =-1114;
9647: waveform_sig_rx =-1288;
9648: waveform_sig_rx =-1135;
9649: waveform_sig_rx =-990;
9650: waveform_sig_rx =-1344;
9651: waveform_sig_rx =-1090;
9652: waveform_sig_rx =-1196;
9653: waveform_sig_rx =-1168;
9654: waveform_sig_rx =-1145;
9655: waveform_sig_rx =-1105;
9656: waveform_sig_rx =-1240;
9657: waveform_sig_rx =-1179;
9658: waveform_sig_rx =-982;
9659: waveform_sig_rx =-1420;
9660: waveform_sig_rx =-1018;
9661: waveform_sig_rx =-1094;
9662: waveform_sig_rx =-1384;
9663: waveform_sig_rx =-1022;
9664: waveform_sig_rx =-1090;
9665: waveform_sig_rx =-1371;
9666: waveform_sig_rx =-1079;
9667: waveform_sig_rx =-1073;
9668: waveform_sig_rx =-1319;
9669: waveform_sig_rx =-1144;
9670: waveform_sig_rx =-1058;
9671: waveform_sig_rx =-1223;
9672: waveform_sig_rx =-1324;
9673: waveform_sig_rx =-963;
9674: waveform_sig_rx =-1196;
9675: waveform_sig_rx =-1300;
9676: waveform_sig_rx =-1077;
9677: waveform_sig_rx =-1071;
9678: waveform_sig_rx =-1361;
9679: waveform_sig_rx =-1093;
9680: waveform_sig_rx =-1075;
9681: waveform_sig_rx =-1247;
9682: waveform_sig_rx =-1188;
9683: waveform_sig_rx =-1044;
9684: waveform_sig_rx =-1150;
9685: waveform_sig_rx =-1310;
9686: waveform_sig_rx =-1024;
9687: waveform_sig_rx =-1108;
9688: waveform_sig_rx =-1339;
9689: waveform_sig_rx =-1060;
9690: waveform_sig_rx =-1024;
9691: waveform_sig_rx =-1345;
9692: waveform_sig_rx =-1022;
9693: waveform_sig_rx =-1237;
9694: waveform_sig_rx =-1126;
9695: waveform_sig_rx =-1148;
9696: waveform_sig_rx =-1111;
9697: waveform_sig_rx =-1240;
9698: waveform_sig_rx =-1138;
9699: waveform_sig_rx =-1008;
9700: waveform_sig_rx =-1380;
9701: waveform_sig_rx =-972;
9702: waveform_sig_rx =-1123;
9703: waveform_sig_rx =-1281;
9704: waveform_sig_rx =-1014;
9705: waveform_sig_rx =-1067;
9706: waveform_sig_rx =-1278;
9707: waveform_sig_rx =-1107;
9708: waveform_sig_rx =-985;
9709: waveform_sig_rx =-1285;
9710: waveform_sig_rx =-1148;
9711: waveform_sig_rx =-944;
9712: waveform_sig_rx =-1236;
9713: waveform_sig_rx =-1220;
9714: waveform_sig_rx =-882;
9715: waveform_sig_rx =-1214;
9716: waveform_sig_rx =-1168;
9717: waveform_sig_rx =-1049;
9718: waveform_sig_rx =-1038;
9719: waveform_sig_rx =-1247;
9720: waveform_sig_rx =-1045;
9721: waveform_sig_rx =-991;
9722: waveform_sig_rx =-1208;
9723: waveform_sig_rx =-1141;
9724: waveform_sig_rx =-965;
9725: waveform_sig_rx =-1101;
9726: waveform_sig_rx =-1245;
9727: waveform_sig_rx =-918;
9728: waveform_sig_rx =-1053;
9729: waveform_sig_rx =-1285;
9730: waveform_sig_rx =-930;
9731: waveform_sig_rx =-1005;
9732: waveform_sig_rx =-1253;
9733: waveform_sig_rx =-914;
9734: waveform_sig_rx =-1209;
9735: waveform_sig_rx =-981;
9736: waveform_sig_rx =-1083;
9737: waveform_sig_rx =-1033;
9738: waveform_sig_rx =-1105;
9739: waveform_sig_rx =-1057;
9740: waveform_sig_rx =-922;
9741: waveform_sig_rx =-1254;
9742: waveform_sig_rx =-931;
9743: waveform_sig_rx =-971;
9744: waveform_sig_rx =-1190;
9745: waveform_sig_rx =-916;
9746: waveform_sig_rx =-909;
9747: waveform_sig_rx =-1247;
9748: waveform_sig_rx =-935;
9749: waveform_sig_rx =-851;
9750: waveform_sig_rx =-1237;
9751: waveform_sig_rx =-955;
9752: waveform_sig_rx =-836;
9753: waveform_sig_rx =-1158;
9754: waveform_sig_rx =-1033;
9755: waveform_sig_rx =-809;
9756: waveform_sig_rx =-1087;
9757: waveform_sig_rx =-1004;
9758: waveform_sig_rx =-942;
9759: waveform_sig_rx =-872;
9760: waveform_sig_rx =-1114;
9761: waveform_sig_rx =-934;
9762: waveform_sig_rx =-833;
9763: waveform_sig_rx =-1076;
9764: waveform_sig_rx =-1006;
9765: waveform_sig_rx =-753;
9766: waveform_sig_rx =-999;
9767: waveform_sig_rx =-1098;
9768: waveform_sig_rx =-716;
9769: waveform_sig_rx =-963;
9770: waveform_sig_rx =-1087;
9771: waveform_sig_rx =-760;
9772: waveform_sig_rx =-900;
9773: waveform_sig_rx =-1026;
9774: waveform_sig_rx =-807;
9775: waveform_sig_rx =-1035;
9776: waveform_sig_rx =-763;
9777: waveform_sig_rx =-982;
9778: waveform_sig_rx =-822;
9779: waveform_sig_rx =-965;
9780: waveform_sig_rx =-922;
9781: waveform_sig_rx =-722;
9782: waveform_sig_rx =-1097;
9783: waveform_sig_rx =-745;
9784: waveform_sig_rx =-776;
9785: waveform_sig_rx =-1085;
9786: waveform_sig_rx =-686;
9787: waveform_sig_rx =-768;
9788: waveform_sig_rx =-1095;
9789: waveform_sig_rx =-693;
9790: waveform_sig_rx =-721;
9791: waveform_sig_rx =-1056;
9792: waveform_sig_rx =-708;
9793: waveform_sig_rx =-697;
9794: waveform_sig_rx =-959;
9795: waveform_sig_rx =-821;
9796: waveform_sig_rx =-662;
9797: waveform_sig_rx =-867;
9798: waveform_sig_rx =-823;
9799: waveform_sig_rx =-785;
9800: waveform_sig_rx =-644;
9801: waveform_sig_rx =-970;
9802: waveform_sig_rx =-731;
9803: waveform_sig_rx =-614;
9804: waveform_sig_rx =-935;
9805: waveform_sig_rx =-767;
9806: waveform_sig_rx =-571;
9807: waveform_sig_rx =-856;
9808: waveform_sig_rx =-804;
9809: waveform_sig_rx =-555;
9810: waveform_sig_rx =-781;
9811: waveform_sig_rx =-814;
9812: waveform_sig_rx =-610;
9813: waveform_sig_rx =-645;
9814: waveform_sig_rx =-811;
9815: waveform_sig_rx =-634;
9816: waveform_sig_rx =-752;
9817: waveform_sig_rx =-592;
9818: waveform_sig_rx =-772;
9819: waveform_sig_rx =-540;
9820: waveform_sig_rx =-788;
9821: waveform_sig_rx =-620;
9822: waveform_sig_rx =-487;
9823: waveform_sig_rx =-918;
9824: waveform_sig_rx =-454;
9825: waveform_sig_rx =-572;
9826: waveform_sig_rx =-850;
9827: waveform_sig_rx =-421;
9828: waveform_sig_rx =-550;
9829: waveform_sig_rx =-861;
9830: waveform_sig_rx =-421;
9831: waveform_sig_rx =-537;
9832: waveform_sig_rx =-805;
9833: waveform_sig_rx =-441;
9834: waveform_sig_rx =-529;
9835: waveform_sig_rx =-673;
9836: waveform_sig_rx =-587;
9837: waveform_sig_rx =-466;
9838: waveform_sig_rx =-571;
9839: waveform_sig_rx =-675;
9840: waveform_sig_rx =-466;
9841: waveform_sig_rx =-390;
9842: waveform_sig_rx =-777;
9843: waveform_sig_rx =-373;
9844: waveform_sig_rx =-423;
9845: waveform_sig_rx =-688;
9846: waveform_sig_rx =-460;
9847: waveform_sig_rx =-384;
9848: waveform_sig_rx =-562;
9849: waveform_sig_rx =-596;
9850: waveform_sig_rx =-338;
9851: waveform_sig_rx =-497;
9852: waveform_sig_rx =-594;
9853: waveform_sig_rx =-356;
9854: waveform_sig_rx =-395;
9855: waveform_sig_rx =-575;
9856: waveform_sig_rx =-376;
9857: waveform_sig_rx =-486;
9858: waveform_sig_rx =-359;
9859: waveform_sig_rx =-487;
9860: waveform_sig_rx =-239;
9861: waveform_sig_rx =-571;
9862: waveform_sig_rx =-314;
9863: waveform_sig_rx =-265;
9864: waveform_sig_rx =-648;
9865: waveform_sig_rx =-126;
9866: waveform_sig_rx =-410;
9867: waveform_sig_rx =-542;
9868: waveform_sig_rx =-114;
9869: waveform_sig_rx =-365;
9870: waveform_sig_rx =-494;
9871: waveform_sig_rx =-188;
9872: waveform_sig_rx =-282;
9873: waveform_sig_rx =-457;
9874: waveform_sig_rx =-240;
9875: waveform_sig_rx =-209;
9876: waveform_sig_rx =-404;
9877: waveform_sig_rx =-352;
9878: waveform_sig_rx =-122;
9879: waveform_sig_rx =-339;
9880: waveform_sig_rx =-371;
9881: waveform_sig_rx =-134;
9882: waveform_sig_rx =-181;
9883: waveform_sig_rx =-452;
9884: waveform_sig_rx =-103;
9885: waveform_sig_rx =-184;
9886: waveform_sig_rx =-370;
9887: waveform_sig_rx =-183;
9888: waveform_sig_rx =-102;
9889: waveform_sig_rx =-267;
9890: waveform_sig_rx =-271;
9891: waveform_sig_rx =-43;
9892: waveform_sig_rx =-174;
9893: waveform_sig_rx =-316;
9894: waveform_sig_rx =-36;
9895: waveform_sig_rx =-60;
9896: waveform_sig_rx =-330;
9897: waveform_sig_rx =-21;
9898: waveform_sig_rx =-196;
9899: waveform_sig_rx =-106;
9900: waveform_sig_rx =-127;
9901: waveform_sig_rx =-29;
9902: waveform_sig_rx =-266;
9903: waveform_sig_rx =48;
9904: waveform_sig_rx =-60;
9905: waveform_sig_rx =-281;
9906: waveform_sig_rx =147;
9907: waveform_sig_rx =-154;
9908: waveform_sig_rx =-177;
9909: waveform_sig_rx =104;
9910: waveform_sig_rx =-35;
9911: waveform_sig_rx =-212;
9912: waveform_sig_rx =64;
9913: waveform_sig_rx =35;
9914: waveform_sig_rx =-208;
9915: waveform_sig_rx =59;
9916: waveform_sig_rx =94;
9917: waveform_sig_rx =-159;
9918: waveform_sig_rx =-21;
9919: waveform_sig_rx =177;
9920: waveform_sig_rx =-66;
9921: waveform_sig_rx =-56;
9922: waveform_sig_rx =147;
9923: waveform_sig_rx =88;
9924: waveform_sig_rx =-122;
9925: waveform_sig_rx =195;
9926: waveform_sig_rx =102;
9927: waveform_sig_rx =-41;
9928: waveform_sig_rx =91;
9929: waveform_sig_rx =208;
9930: waveform_sig_rx =31;
9931: waveform_sig_rx =-18;
9932: waveform_sig_rx =290;
9933: waveform_sig_rx =95;
9934: waveform_sig_rx =-76;
9935: waveform_sig_rx =311;
9936: waveform_sig_rx =156;
9937: waveform_sig_rx =-34;
9938: waveform_sig_rx =316;
9939: waveform_sig_rx =-4;
9940: waveform_sig_rx =266;
9941: waveform_sig_rx =144;
9942: waveform_sig_rx =226;
9943: waveform_sig_rx =94;
9944: waveform_sig_rx =280;
9945: waveform_sig_rx =222;
9946: waveform_sig_rx =35;
9947: waveform_sig_rx =350;
9948: waveform_sig_rx =205;
9949: waveform_sig_rx =44;
9950: waveform_sig_rx =400;
9951: waveform_sig_rx =267;
9952: waveform_sig_rx =20;
9953: waveform_sig_rx =448;
9954: waveform_sig_rx =280;
9955: waveform_sig_rx =99;
9956: waveform_sig_rx =359;
9957: waveform_sig_rx =391;
9958: waveform_sig_rx =127;
9959: waveform_sig_rx =270;
9960: waveform_sig_rx =522;
9961: waveform_sig_rx =152;
9962: waveform_sig_rx =281;
9963: waveform_sig_rx =445;
9964: waveform_sig_rx =315;
9965: waveform_sig_rx =248;
9966: waveform_sig_rx =399;
9967: waveform_sig_rx =439;
9968: waveform_sig_rx =249;
9969: waveform_sig_rx =318;
9970: waveform_sig_rx =607;
9971: waveform_sig_rx =234;
9972: waveform_sig_rx =297;
9973: waveform_sig_rx =623;
9974: waveform_sig_rx =283;
9975: waveform_sig_rx =320;
9976: waveform_sig_rx =567;
9977: waveform_sig_rx =397;
9978: waveform_sig_rx =326;
9979: waveform_sig_rx =510;
9980: waveform_sig_rx =324;
9981: waveform_sig_rx =571;
9982: waveform_sig_rx =381;
9983: waveform_sig_rx =546;
9984: waveform_sig_rx =355;
9985: waveform_sig_rx =539;
9986: waveform_sig_rx =549;
9987: waveform_sig_rx =312;
9988: waveform_sig_rx =658;
9989: waveform_sig_rx =518;
9990: waveform_sig_rx =313;
9991: waveform_sig_rx =714;
9992: waveform_sig_rx =549;
9993: waveform_sig_rx =293;
9994: waveform_sig_rx =746;
9995: waveform_sig_rx =564;
9996: waveform_sig_rx =347;
9997: waveform_sig_rx =698;
9998: waveform_sig_rx =645;
9999: waveform_sig_rx =373;
10000: waveform_sig_rx =610;
10001: waveform_sig_rx =709;
10002: waveform_sig_rx =459;
10003: waveform_sig_rx =585;
10004: waveform_sig_rx =658;
10005: waveform_sig_rx =673;
10006: waveform_sig_rx =448;
10007: waveform_sig_rx =701;
10008: waveform_sig_rx =780;
10009: waveform_sig_rx =438;
10010: waveform_sig_rx =680;
10011: waveform_sig_rx =840;
10012: waveform_sig_rx =438;
10013: waveform_sig_rx =663;
10014: waveform_sig_rx =813;
10015: waveform_sig_rx =574;
10016: waveform_sig_rx =602;
10017: waveform_sig_rx =795;
10018: waveform_sig_rx =721;
10019: waveform_sig_rx =570;
10020: waveform_sig_rx =783;
10021: waveform_sig_rx =617;
10022: waveform_sig_rx =781;
10023: waveform_sig_rx =619;
10024: waveform_sig_rx =815;
10025: waveform_sig_rx =575;
10026: waveform_sig_rx =819;
10027: waveform_sig_rx =768;
10028: waveform_sig_rx =537;
10029: waveform_sig_rx =928;
10030: waveform_sig_rx =736;
10031: waveform_sig_rx =536;
10032: waveform_sig_rx =999;
10033: waveform_sig_rx =754;
10034: waveform_sig_rx =525;
10035: waveform_sig_rx =1045;
10036: waveform_sig_rx =713;
10037: waveform_sig_rx =629;
10038: waveform_sig_rx =947;
10039: waveform_sig_rx =797;
10040: waveform_sig_rx =670;
10041: waveform_sig_rx =819;
10042: waveform_sig_rx =924;
10043: waveform_sig_rx =749;
10044: waveform_sig_rx =738;
10045: waveform_sig_rx =937;
10046: waveform_sig_rx =895;
10047: waveform_sig_rx =618;
10048: waveform_sig_rx =1006;
10049: waveform_sig_rx =891;
10050: waveform_sig_rx =660;
10051: waveform_sig_rx =946;
10052: waveform_sig_rx =978;
10053: waveform_sig_rx =704;
10054: waveform_sig_rx =874;
10055: waveform_sig_rx =1004;
10056: waveform_sig_rx =801;
10057: waveform_sig_rx =789;
10058: waveform_sig_rx =1005;
10059: waveform_sig_rx =899;
10060: waveform_sig_rx =768;
10061: waveform_sig_rx =960;
10062: waveform_sig_rx =836;
10063: waveform_sig_rx =967;
10064: waveform_sig_rx =834;
10065: waveform_sig_rx =1039;
10066: waveform_sig_rx =718;
10067: waveform_sig_rx =1071;
10068: waveform_sig_rx =930;
10069: waveform_sig_rx =708;
10070: waveform_sig_rx =1176;
10071: waveform_sig_rx =841;
10072: waveform_sig_rx =770;
10073: waveform_sig_rx =1226;
10074: waveform_sig_rx =830;
10075: waveform_sig_rx =794;
10076: waveform_sig_rx =1190;
10077: waveform_sig_rx =875;
10078: waveform_sig_rx =897;
10079: waveform_sig_rx =1067;
10080: waveform_sig_rx =1036;
10081: waveform_sig_rx =856;
10082: waveform_sig_rx =975;
10083: waveform_sig_rx =1166;
10084: waveform_sig_rx =886;
10085: waveform_sig_rx =903;
10086: waveform_sig_rx =1162;
10087: waveform_sig_rx =991;
10088: waveform_sig_rx =814;
10089: waveform_sig_rx =1195;
10090: waveform_sig_rx =1010;
10091: waveform_sig_rx =846;
10092: waveform_sig_rx =1128;
10093: waveform_sig_rx =1088;
10094: waveform_sig_rx =894;
10095: waveform_sig_rx =995;
10096: waveform_sig_rx =1149;
10097: waveform_sig_rx =979;
10098: waveform_sig_rx =889;
10099: waveform_sig_rx =1191;
10100: waveform_sig_rx =1035;
10101: waveform_sig_rx =891;
10102: waveform_sig_rx =1176;
10103: waveform_sig_rx =964;
10104: waveform_sig_rx =1118;
10105: waveform_sig_rx =1031;
10106: waveform_sig_rx =1142;
10107: waveform_sig_rx =873;
10108: waveform_sig_rx =1282;
10109: waveform_sig_rx =1021;
10110: waveform_sig_rx =938;
10111: waveform_sig_rx =1330;
10112: waveform_sig_rx =930;
10113: waveform_sig_rx =992;
10114: waveform_sig_rx =1316;
10115: waveform_sig_rx =970;
10116: waveform_sig_rx =990;
10117: waveform_sig_rx =1275;
10118: waveform_sig_rx =1032;
10119: waveform_sig_rx =1008;
10120: waveform_sig_rx =1159;
10121: waveform_sig_rx =1199;
10122: waveform_sig_rx =908;
10123: waveform_sig_rx =1103;
10124: waveform_sig_rx =1277;
10125: waveform_sig_rx =930;
10126: waveform_sig_rx =1078;
10127: waveform_sig_rx =1258;
10128: waveform_sig_rx =1048;
10129: waveform_sig_rx =995;
10130: waveform_sig_rx =1265;
10131: waveform_sig_rx =1097;
10132: waveform_sig_rx =984;
10133: waveform_sig_rx =1177;
10134: waveform_sig_rx =1224;
10135: waveform_sig_rx =995;
10136: waveform_sig_rx =1086;
10137: waveform_sig_rx =1281;
10138: waveform_sig_rx =1045;
10139: waveform_sig_rx =1004;
10140: waveform_sig_rx =1345;
10141: waveform_sig_rx =1089;
10142: waveform_sig_rx =1026;
10143: waveform_sig_rx =1278;
10144: waveform_sig_rx =997;
10145: waveform_sig_rx =1230;
10146: waveform_sig_rx =1115;
10147: waveform_sig_rx =1187;
10148: waveform_sig_rx =1002;
10149: waveform_sig_rx =1352;
10150: waveform_sig_rx =1040;
10151: waveform_sig_rx =1062;
10152: waveform_sig_rx =1332;
10153: waveform_sig_rx =1010;
10154: waveform_sig_rx =1098;
10155: waveform_sig_rx =1316;
10156: waveform_sig_rx =1086;
10157: waveform_sig_rx =1017;
10158: waveform_sig_rx =1321;
10159: waveform_sig_rx =1133;
10160: waveform_sig_rx =999;
10161: waveform_sig_rx =1264;
10162: waveform_sig_rx =1230;
10163: waveform_sig_rx =907;
10164: waveform_sig_rx =1254;
10165: waveform_sig_rx =1245;
10166: waveform_sig_rx =988;
10167: waveform_sig_rx =1148;
10168: waveform_sig_rx =1242;
10169: waveform_sig_rx =1120;
10170: waveform_sig_rx =1029;
10171: waveform_sig_rx =1285;
10172: waveform_sig_rx =1166;
10173: waveform_sig_rx =1020;
10174: waveform_sig_rx =1205;
10175: waveform_sig_rx =1285;
10176: waveform_sig_rx =1003;
10177: waveform_sig_rx =1137;
10178: waveform_sig_rx =1341;
10179: waveform_sig_rx =1025;
10180: waveform_sig_rx =1060;
10181: waveform_sig_rx =1373;
10182: waveform_sig_rx =1032;
10183: waveform_sig_rx =1102;
10184: waveform_sig_rx =1251;
10185: waveform_sig_rx =1002;
10186: waveform_sig_rx =1272;
10187: waveform_sig_rx =1052;
10188: waveform_sig_rx =1205;
10189: waveform_sig_rx =1006;
10190: waveform_sig_rx =1295;
10191: waveform_sig_rx =1057;
10192: waveform_sig_rx =1043;
10193: waveform_sig_rx =1296;
10194: waveform_sig_rx =1062;
10195: waveform_sig_rx =1021;
10196: waveform_sig_rx =1336;
10197: waveform_sig_rx =1072;
10198: waveform_sig_rx =936;
10199: waveform_sig_rx =1381;
10200: waveform_sig_rx =1045;
10201: waveform_sig_rx =977;
10202: waveform_sig_rx =1309;
10203: waveform_sig_rx =1133;
10204: waveform_sig_rx =942;
10205: waveform_sig_rx =1242;
10206: waveform_sig_rx =1174;
10207: waveform_sig_rx =1026;
10208: waveform_sig_rx =1083;
10209: waveform_sig_rx =1230;
10210: waveform_sig_rx =1068;
10211: waveform_sig_rx =966;
10212: waveform_sig_rx =1283;
10213: waveform_sig_rx =1100;
10214: waveform_sig_rx =972;
10215: waveform_sig_rx =1154;
10216: waveform_sig_rx =1238;
10217: waveform_sig_rx =885;
10218: waveform_sig_rx =1093;
10219: waveform_sig_rx =1296;
10220: waveform_sig_rx =893;
10221: waveform_sig_rx =1089;
10222: waveform_sig_rx =1246;
10223: waveform_sig_rx =961;
10224: waveform_sig_rx =1116;
10225: waveform_sig_rx =1051;
10226: waveform_sig_rx =1035;
10227: waveform_sig_rx =1181;
10228: waveform_sig_rx =949;
10229: waveform_sig_rx =1215;
10230: waveform_sig_rx =869;
10231: waveform_sig_rx =1255;
10232: waveform_sig_rx =1011;
10233: waveform_sig_rx =898;
10234: waveform_sig_rx =1284;
10235: waveform_sig_rx =925;
10236: waveform_sig_rx =945;
10237: waveform_sig_rx =1281;
10238: waveform_sig_rx =921;
10239: waveform_sig_rx =894;
10240: waveform_sig_rx =1277;
10241: waveform_sig_rx =924;
10242: waveform_sig_rx =900;
10243: waveform_sig_rx =1216;
10244: waveform_sig_rx =984;
10245: waveform_sig_rx =840;
10246: waveform_sig_rx =1136;
10247: waveform_sig_rx =1026;
10248: waveform_sig_rx =956;
10249: waveform_sig_rx =940;
10250: waveform_sig_rx =1133;
10251: waveform_sig_rx =976;
10252: waveform_sig_rx =827;
10253: waveform_sig_rx =1187;
10254: waveform_sig_rx =961;
10255: waveform_sig_rx =820;
10256: waveform_sig_rx =1117;
10257: waveform_sig_rx =1052;
10258: waveform_sig_rx =784;
10259: waveform_sig_rx =1058;
10260: waveform_sig_rx =1092;
10261: waveform_sig_rx =825;
10262: waveform_sig_rx =949;
10263: waveform_sig_rx =1075;
10264: waveform_sig_rx =895;
10265: waveform_sig_rx =912;
10266: waveform_sig_rx =938;
10267: waveform_sig_rx =936;
10268: waveform_sig_rx =969;
10269: waveform_sig_rx =890;
10270: waveform_sig_rx =1047;
10271: waveform_sig_rx =688;
10272: waveform_sig_rx =1164;
10273: waveform_sig_rx =785;
10274: waveform_sig_rx =795;
10275: waveform_sig_rx =1157;
10276: waveform_sig_rx =710;
10277: waveform_sig_rx =856;
10278: waveform_sig_rx =1102;
10279: waveform_sig_rx =743;
10280: waveform_sig_rx =767;
10281: waveform_sig_rx =1113;
10282: waveform_sig_rx =734;
10283: waveform_sig_rx =787;
10284: waveform_sig_rx =1036;
10285: waveform_sig_rx =832;
10286: waveform_sig_rx =735;
10287: waveform_sig_rx =955;
10288: waveform_sig_rx =898;
10289: waveform_sig_rx =789;
10290: waveform_sig_rx =726;
10291: waveform_sig_rx =1023;
10292: waveform_sig_rx =756;
10293: waveform_sig_rx =676;
10294: waveform_sig_rx =1064;
10295: waveform_sig_rx =706;
10296: waveform_sig_rx =700;
10297: waveform_sig_rx =916;
10298: waveform_sig_rx =812;
10299: waveform_sig_rx =668;
10300: waveform_sig_rx =785;
10301: waveform_sig_rx =884;
10302: waveform_sig_rx =658;
10303: waveform_sig_rx =703;
10304: waveform_sig_rx =944;
10305: waveform_sig_rx =650;
10306: waveform_sig_rx =698;
10307: waveform_sig_rx =780;
10308: waveform_sig_rx =687;
10309: waveform_sig_rx =765;
10310: waveform_sig_rx =691;
10311: waveform_sig_rx =779;
10312: waveform_sig_rx =531;
10313: waveform_sig_rx =959;
10314: waveform_sig_rx =540;
10315: waveform_sig_rx =656;
10316: waveform_sig_rx =930;
10317: waveform_sig_rx =471;
10318: waveform_sig_rx =681;
10319: waveform_sig_rx =873;
10320: waveform_sig_rx =496;
10321: waveform_sig_rx =630;
10322: waveform_sig_rx =845;
10323: waveform_sig_rx =528;
10324: waveform_sig_rx =623;
10325: waveform_sig_rx =731;
10326: waveform_sig_rx =665;
10327: waveform_sig_rx =453;
10328: waveform_sig_rx =696;
10329: waveform_sig_rx =705;
10330: waveform_sig_rx =443;
10331: waveform_sig_rx =562;
10332: waveform_sig_rx =772;
10333: waveform_sig_rx =439;
10334: waveform_sig_rx =512;
10335: waveform_sig_rx =734;
10336: waveform_sig_rx =491;
10337: waveform_sig_rx =483;
10338: waveform_sig_rx =635;
10339: waveform_sig_rx =610;
10340: waveform_sig_rx =389;
10341: waveform_sig_rx =552;
10342: waveform_sig_rx =648;
10343: waveform_sig_rx =394;
10344: waveform_sig_rx =446;
10345: waveform_sig_rx =716;
10346: waveform_sig_rx =389;
10347: waveform_sig_rx =458;
10348: waveform_sig_rx =570;
10349: waveform_sig_rx =398;
10350: waveform_sig_rx =520;
10351: waveform_sig_rx =464;
10352: waveform_sig_rx =467;
10353: waveform_sig_rx =319;
10354: waveform_sig_rx =691;
10355: waveform_sig_rx =232;
10356: waveform_sig_rx =441;
10357: waveform_sig_rx =587;
10358: waveform_sig_rx =246;
10359: waveform_sig_rx =435;
10360: waveform_sig_rx =551;
10361: waveform_sig_rx =281;
10362: waveform_sig_rx =320;
10363: waveform_sig_rx =569;
10364: waveform_sig_rx =303;
10365: waveform_sig_rx =284;
10366: waveform_sig_rx =501;
10367: waveform_sig_rx =379;
10368: waveform_sig_rx =151;
10369: waveform_sig_rx =490;
10370: waveform_sig_rx =387;
10371: waveform_sig_rx =180;
10372: waveform_sig_rx =351;
10373: waveform_sig_rx =453;
10374: waveform_sig_rx =190;
10375: waveform_sig_rx =276;
10376: waveform_sig_rx =442;
10377: waveform_sig_rx =234;
10378: waveform_sig_rx =196;
10379: waveform_sig_rx =349;
10380: waveform_sig_rx =354;
10381: waveform_sig_rx =84;
10382: waveform_sig_rx =288;
10383: waveform_sig_rx =410;
10384: waveform_sig_rx =56;
10385: waveform_sig_rx =198;
10386: waveform_sig_rx =412;
10387: waveform_sig_rx =14;
10388: waveform_sig_rx =234;
10389: waveform_sig_rx =213;
10390: waveform_sig_rx =107;
10391: waveform_sig_rx =283;
10392: waveform_sig_rx =131;
10393: waveform_sig_rx =198;
10394: waveform_sig_rx =53;
10395: waveform_sig_rx =333;
10396: waveform_sig_rx =-10;
10397: waveform_sig_rx =137;
10398: waveform_sig_rx =262;
10399: waveform_sig_rx =-11;
10400: waveform_sig_rx =89;
10401: waveform_sig_rx =292;
10402: waveform_sig_rx =-44;
10403: waveform_sig_rx =3;
10404: waveform_sig_rx =320;
10405: waveform_sig_rx =-72;
10406: waveform_sig_rx =-4;
10407: waveform_sig_rx =211;
10408: waveform_sig_rx =28;
10409: waveform_sig_rx =-146;
10410: waveform_sig_rx =218;
10411: waveform_sig_rx =40;
10412: waveform_sig_rx =-107;
10413: waveform_sig_rx =53;
10414: waveform_sig_rx =113;
10415: waveform_sig_rx =-97;
10416: waveform_sig_rx =-68;
10417: waveform_sig_rx =108;
10418: waveform_sig_rx =-45;
10419: waveform_sig_rx =-185;
10420: waveform_sig_rx =71;
10421: waveform_sig_rx =58;
10422: waveform_sig_rx =-309;
10423: waveform_sig_rx =58;
10424: waveform_sig_rx =47;
10425: waveform_sig_rx =-281;
10426: waveform_sig_rx =-32;
10427: waveform_sig_rx =30;
10428: waveform_sig_rx =-242;
10429: waveform_sig_rx =-53;
10430: waveform_sig_rx =-154;
10431: waveform_sig_rx =-122;
10432: waveform_sig_rx =-75;
10433: waveform_sig_rx =-180;
10434: waveform_sig_rx =-67;
10435: waveform_sig_rx =-289;
10436: waveform_sig_rx =35;
10437: waveform_sig_rx =-287;
10438: waveform_sig_rx =-194;
10439: waveform_sig_rx =19;
10440: waveform_sig_rx =-349;
10441: waveform_sig_rx =-215;
10442: waveform_sig_rx =14;
10443: waveform_sig_rx =-392;
10444: waveform_sig_rx =-290;
10445: waveform_sig_rx =13;
10446: waveform_sig_rx =-416;
10447: waveform_sig_rx =-293;
10448: waveform_sig_rx =-69;
10449: waveform_sig_rx =-321;
10450: waveform_sig_rx =-420;
10451: waveform_sig_rx =-92;
10452: waveform_sig_rx =-319;
10453: waveform_sig_rx =-360;
10454: waveform_sig_rx =-295;
10455: waveform_sig_rx =-173;
10456: waveform_sig_rx =-363;
10457: waveform_sig_rx =-433;
10458: waveform_sig_rx =-136;
10459: waveform_sig_rx =-387;
10460: waveform_sig_rx =-509;
10461: waveform_sig_rx =-147;
10462: waveform_sig_rx =-364;
10463: waveform_sig_rx =-550;
10464: waveform_sig_rx =-219;
10465: waveform_sig_rx =-339;
10466: waveform_sig_rx =-495;
10467: waveform_sig_rx =-384;
10468: waveform_sig_rx =-250;
10469: waveform_sig_rx =-511;
10470: waveform_sig_rx =-399;
10471: waveform_sig_rx =-428;
10472: waveform_sig_rx =-427;
10473: waveform_sig_rx =-398;
10474: waveform_sig_rx =-455;
10475: waveform_sig_rx =-380;
10476: waveform_sig_rx =-612;
10477: waveform_sig_rx =-249;
10478: waveform_sig_rx =-637;
10479: waveform_sig_rx =-522;
10480: waveform_sig_rx =-261;
10481: waveform_sig_rx =-707;
10482: waveform_sig_rx =-518;
10483: waveform_sig_rx =-235;
10484: waveform_sig_rx =-777;
10485: waveform_sig_rx =-501;
10486: waveform_sig_rx =-287;
10487: waveform_sig_rx =-765;
10488: waveform_sig_rx =-482;
10489: waveform_sig_rx =-450;
10490: waveform_sig_rx =-567;
10491: waveform_sig_rx =-665;
10492: waveform_sig_rx =-443;
10493: waveform_sig_rx =-536;
10494: waveform_sig_rx =-678;
10495: waveform_sig_rx =-596;
10496: waveform_sig_rx =-414;
10497: waveform_sig_rx =-725;
10498: waveform_sig_rx =-683;
10499: waveform_sig_rx =-399;
10500: waveform_sig_rx =-724;
10501: waveform_sig_rx =-736;
10502: waveform_sig_rx =-433;
10503: waveform_sig_rx =-657;
10504: waveform_sig_rx =-768;
10505: waveform_sig_rx =-529;
10506: waveform_sig_rx =-617;
10507: waveform_sig_rx =-759;
10508: waveform_sig_rx =-697;
10509: waveform_sig_rx =-494;
10510: waveform_sig_rx =-800;
10511: waveform_sig_rx =-685;
10512: waveform_sig_rx =-665;
10513: waveform_sig_rx =-695;
10514: waveform_sig_rx =-705;
10515: waveform_sig_rx =-691;
10516: waveform_sig_rx =-710;
10517: waveform_sig_rx =-847;
10518: waveform_sig_rx =-474;
10519: waveform_sig_rx =-941;
10520: waveform_sig_rx =-718;
10521: waveform_sig_rx =-538;
10522: waveform_sig_rx =-1019;
10523: waveform_sig_rx =-676;
10524: waveform_sig_rx =-575;
10525: waveform_sig_rx =-1041;
10526: waveform_sig_rx =-683;
10527: waveform_sig_rx =-641;
10528: waveform_sig_rx =-970;
10529: waveform_sig_rx =-744;
10530: waveform_sig_rx =-730;
10531: waveform_sig_rx =-768;
10532: waveform_sig_rx =-984;
10533: waveform_sig_rx =-667;
10534: waveform_sig_rx =-774;
10535: waveform_sig_rx =-982;
10536: waveform_sig_rx =-790;
10537: waveform_sig_rx =-692;
10538: waveform_sig_rx =-1030;
10539: waveform_sig_rx =-859;
10540: waveform_sig_rx =-673;
10541: waveform_sig_rx =-972;
10542: waveform_sig_rx =-932;
10543: waveform_sig_rx =-709;
10544: waveform_sig_rx =-889;
10545: waveform_sig_rx =-979;
10546: waveform_sig_rx =-772;
10547: waveform_sig_rx =-810;
10548: waveform_sig_rx =-990;
10549: waveform_sig_rx =-925;
10550: waveform_sig_rx =-689;
10551: waveform_sig_rx =-1063;
10552: waveform_sig_rx =-889;
10553: waveform_sig_rx =-873;
10554: waveform_sig_rx =-962;
10555: waveform_sig_rx =-885;
10556: waveform_sig_rx =-888;
10557: waveform_sig_rx =-995;
10558: waveform_sig_rx =-1000;
10559: waveform_sig_rx =-737;
10560: waveform_sig_rx =-1196;
10561: waveform_sig_rx =-857;
10562: waveform_sig_rx =-836;
10563: waveform_sig_rx =-1170;
10564: waveform_sig_rx =-861;
10565: waveform_sig_rx =-844;
10566: waveform_sig_rx =-1158;
10567: waveform_sig_rx =-920;
10568: waveform_sig_rx =-848;
10569: waveform_sig_rx =-1130;
10570: waveform_sig_rx =-990;
10571: waveform_sig_rx =-872;
10572: waveform_sig_rx =-994;
10573: waveform_sig_rx =-1184;
10574: waveform_sig_rx =-810;
10575: waveform_sig_rx =-1012;
10576: waveform_sig_rx =-1167;
10577: waveform_sig_rx =-924;
10578: waveform_sig_rx =-908;
10579: waveform_sig_rx =-1192;
10580: waveform_sig_rx =-1004;
10581: waveform_sig_rx =-925;
10582: waveform_sig_rx =-1148;
10583: waveform_sig_rx =-1103;
10584: waveform_sig_rx =-946;
10585: waveform_sig_rx =-1018;
10586: waveform_sig_rx =-1222;
10587: waveform_sig_rx =-966;
10588: waveform_sig_rx =-968;
10589: waveform_sig_rx =-1264;
10590: waveform_sig_rx =-1019;
10591: waveform_sig_rx =-895;
10592: waveform_sig_rx =-1277;
10593: waveform_sig_rx =-983;
10594: waveform_sig_rx =-1108;
10595: waveform_sig_rx =-1094;
10596: waveform_sig_rx =-1037;
10597: waveform_sig_rx =-1087;
10598: waveform_sig_rx =-1116;
10599: waveform_sig_rx =-1123;
10600: waveform_sig_rx =-932;
10601: waveform_sig_rx =-1315;
10602: waveform_sig_rx =-1023;
10603: waveform_sig_rx =-1041;
10604: waveform_sig_rx =-1282;
10605: waveform_sig_rx =-1028;
10606: waveform_sig_rx =-999;
10607: waveform_sig_rx =-1280;
10608: waveform_sig_rx =-1123;
10609: waveform_sig_rx =-922;
10610: waveform_sig_rx =-1274;
10611: waveform_sig_rx =-1155;
10612: waveform_sig_rx =-937;
10613: waveform_sig_rx =-1204;
10614: waveform_sig_rx =-1298;
10615: waveform_sig_rx =-901;
10616: waveform_sig_rx =-1200;
10617: waveform_sig_rx =-1206;
10618: waveform_sig_rx =-1081;
10619: waveform_sig_rx =-1050;
10620: waveform_sig_rx =-1267;
10621: waveform_sig_rx =-1132;
10622: waveform_sig_rx =-1005;
10623: waveform_sig_rx =-1230;
10624: waveform_sig_rx =-1230;
10625: waveform_sig_rx =-1001;
10626: waveform_sig_rx =-1123;
10627: waveform_sig_rx =-1338;
10628: waveform_sig_rx =-1010;
10629: waveform_sig_rx =-1093;
10630: waveform_sig_rx =-1375;
10631: waveform_sig_rx =-1056;
10632: waveform_sig_rx =-1040;
10633: waveform_sig_rx =-1358;
10634: waveform_sig_rx =-1010;
10635: waveform_sig_rx =-1269;
10636: waveform_sig_rx =-1127;
10637: waveform_sig_rx =-1140;
10638: waveform_sig_rx =-1192;
10639: waveform_sig_rx =-1176;
10640: waveform_sig_rx =-1244;
10641: waveform_sig_rx =-1014;
10642: waveform_sig_rx =-1351;
10643: waveform_sig_rx =-1114;
10644: waveform_sig_rx =-1050;
10645: waveform_sig_rx =-1341;
10646: waveform_sig_rx =-1118;
10647: waveform_sig_rx =-983;
10648: waveform_sig_rx =-1366;
10649: waveform_sig_rx =-1132;
10650: waveform_sig_rx =-947;
10651: waveform_sig_rx =-1422;
10652: waveform_sig_rx =-1129;
10653: waveform_sig_rx =-985;
10654: waveform_sig_rx =-1323;
10655: waveform_sig_rx =-1242;
10656: waveform_sig_rx =-989;
10657: waveform_sig_rx =-1245;
10658: waveform_sig_rx =-1212;
10659: waveform_sig_rx =-1156;
10660: waveform_sig_rx =-1041;
10661: waveform_sig_rx =-1300;
10662: waveform_sig_rx =-1177;
10663: waveform_sig_rx =-1001;
10664: waveform_sig_rx =-1276;
10665: waveform_sig_rx =-1245;
10666: waveform_sig_rx =-994;
10667: waveform_sig_rx =-1187;
10668: waveform_sig_rx =-1347;
10669: waveform_sig_rx =-980;
10670: waveform_sig_rx =-1150;
10671: waveform_sig_rx =-1347;
10672: waveform_sig_rx =-1030;
10673: waveform_sig_rx =-1109;
10674: waveform_sig_rx =-1295;
10675: waveform_sig_rx =-1062;
10676: waveform_sig_rx =-1286;
10677: waveform_sig_rx =-1033;
10678: waveform_sig_rx =-1213;
10679: waveform_sig_rx =-1121;
10680: waveform_sig_rx =-1137;
10681: waveform_sig_rx =-1266;
10682: waveform_sig_rx =-924;
10683: waveform_sig_rx =-1357;
10684: waveform_sig_rx =-1092;
10685: waveform_sig_rx =-977;
10686: waveform_sig_rx =-1402;
10687: waveform_sig_rx =-1020;
10688: waveform_sig_rx =-991;
10689: waveform_sig_rx =-1400;
10690: waveform_sig_rx =-1026;
10691: waveform_sig_rx =-992;
10692: waveform_sig_rx =-1357;
10693: waveform_sig_rx =-1057;
10694: waveform_sig_rx =-1004;
10695: waveform_sig_rx =-1249;
10696: waveform_sig_rx =-1195;
10697: waveform_sig_rx =-966;
10698: waveform_sig_rx =-1168;
10699: waveform_sig_rx =-1181;
10700: waveform_sig_rx =-1104;
10701: waveform_sig_rx =-947;
10702: waveform_sig_rx =-1275;
10703: waveform_sig_rx =-1099;
10704: waveform_sig_rx =-901;
10705: waveform_sig_rx =-1254;
10706: waveform_sig_rx =-1153;
10707: waveform_sig_rx =-881;
10708: waveform_sig_rx =-1182;
10709: waveform_sig_rx =-1197;
10710: waveform_sig_rx =-898;
10711: waveform_sig_rx =-1116;
10712: waveform_sig_rx =-1158;
10713: waveform_sig_rx =-1020;
10714: waveform_sig_rx =-968;
10715: waveform_sig_rx =-1174;
10716: waveform_sig_rx =-1050;
10717: waveform_sig_rx =-1085;
10718: waveform_sig_rx =-984;
10719: waveform_sig_rx =-1141;
10720: waveform_sig_rx =-916;
10721: waveform_sig_rx =-1144;
10722: waveform_sig_rx =-1074;
10723: waveform_sig_rx =-823;
10724: waveform_sig_rx =-1327;
10725: waveform_sig_rx =-879;
10726: waveform_sig_rx =-957;
10727: waveform_sig_rx =-1268;
10728: waveform_sig_rx =-871;
10729: waveform_sig_rx =-920;
10730: waveform_sig_rx =-1249;
10731: waveform_sig_rx =-899;
10732: waveform_sig_rx =-877;
10733: waveform_sig_rx =-1231;
10734: waveform_sig_rx =-900;
10735: waveform_sig_rx =-923;
10736: waveform_sig_rx =-1094;
10737: waveform_sig_rx =-1038;
10738: waveform_sig_rx =-887;
10739: waveform_sig_rx =-974;
10740: waveform_sig_rx =-1073;
10741: waveform_sig_rx =-939;
10742: waveform_sig_rx =-764;
10743: waveform_sig_rx =-1216;
10744: waveform_sig_rx =-855;
10745: waveform_sig_rx =-824;
10746: waveform_sig_rx =-1152;
10747: waveform_sig_rx =-895;
10748: waveform_sig_rx =-862;
10749: waveform_sig_rx =-1001;
10750: waveform_sig_rx =-1031;
10751: waveform_sig_rx =-834;
10752: waveform_sig_rx =-878;
10753: waveform_sig_rx =-1066;
10754: waveform_sig_rx =-858;
10755: waveform_sig_rx =-785;
10756: waveform_sig_rx =-1072;
10757: waveform_sig_rx =-796;
10758: waveform_sig_rx =-954;
10759: waveform_sig_rx =-846;
10760: waveform_sig_rx =-920;
10761: waveform_sig_rx =-791;
10762: waveform_sig_rx =-1017;
10763: waveform_sig_rx =-859;
10764: waveform_sig_rx =-732;
10765: waveform_sig_rx =-1129;
10766: waveform_sig_rx =-674;
10767: waveform_sig_rx =-814;
10768: waveform_sig_rx =-1065;
10769: waveform_sig_rx =-657;
10770: waveform_sig_rx =-789;
10771: waveform_sig_rx =-1029;
10772: waveform_sig_rx =-673;
10773: waveform_sig_rx =-761;
10774: waveform_sig_rx =-985;
10775: waveform_sig_rx =-739;
10776: waveform_sig_rx =-736;
10777: waveform_sig_rx =-850;
10778: waveform_sig_rx =-905;
10779: waveform_sig_rx =-630;
10780: waveform_sig_rx =-792;
10781: waveform_sig_rx =-933;
10782: waveform_sig_rx =-667;
10783: waveform_sig_rx =-674;
10784: waveform_sig_rx =-1015;
10785: waveform_sig_rx =-617;
10786: waveform_sig_rx =-709;
10787: waveform_sig_rx =-887;
10788: waveform_sig_rx =-739;
10789: waveform_sig_rx =-664;
10790: waveform_sig_rx =-733;
10791: waveform_sig_rx =-879;
10792: waveform_sig_rx =-565;
10793: waveform_sig_rx =-674;
10794: waveform_sig_rx =-908;
10795: waveform_sig_rx =-577;
10796: waveform_sig_rx =-617;
10797: waveform_sig_rx =-861;
10798: waveform_sig_rx =-568;
10799: waveform_sig_rx =-770;
10800: waveform_sig_rx =-630;
10801: waveform_sig_rx =-696;
10802: waveform_sig_rx =-581;
10803: waveform_sig_rx =-777;
10804: waveform_sig_rx =-574;
10805: waveform_sig_rx =-541;
10806: waveform_sig_rx =-873;
10807: waveform_sig_rx =-439;
10808: waveform_sig_rx =-642;
10809: waveform_sig_rx =-775;
10810: waveform_sig_rx =-467;
10811: waveform_sig_rx =-582;
10812: waveform_sig_rx =-757;
10813: waveform_sig_rx =-516;
10814: waveform_sig_rx =-461;
10815: waveform_sig_rx =-741;
10816: waveform_sig_rx =-544;
10817: waveform_sig_rx =-405;
10818: waveform_sig_rx =-696;
10819: waveform_sig_rx =-643;
10820: waveform_sig_rx =-336;
10821: waveform_sig_rx =-638;
10822: waveform_sig_rx =-611;
10823: waveform_sig_rx =-427;
10824: waveform_sig_rx =-478;
10825: waveform_sig_rx =-693;
10826: waveform_sig_rx =-447;
10827: waveform_sig_rx =-437;
10828: waveform_sig_rx =-604;
10829: waveform_sig_rx =-526;
10830: waveform_sig_rx =-346;
10831: waveform_sig_rx =-512;
10832: waveform_sig_rx =-633;
10833: waveform_sig_rx =-297;
10834: waveform_sig_rx =-452;
10835: waveform_sig_rx =-654;
10836: waveform_sig_rx =-292;
10837: waveform_sig_rx =-357;
10838: waveform_sig_rx =-627;
10839: waveform_sig_rx =-268;
10840: waveform_sig_rx =-551;
10841: waveform_sig_rx =-344;
10842: waveform_sig_rx =-426;
10843: waveform_sig_rx =-353;
10844: waveform_sig_rx =-488;
10845: waveform_sig_rx =-345;
10846: waveform_sig_rx =-301;
10847: waveform_sig_rx =-551;
10848: waveform_sig_rx =-229;
10849: waveform_sig_rx =-344;
10850: waveform_sig_rx =-506;
10851: waveform_sig_rx =-231;
10852: waveform_sig_rx =-249;
10853: waveform_sig_rx =-544;
10854: waveform_sig_rx =-204;
10855: waveform_sig_rx =-198;
10856: waveform_sig_rx =-524;
10857: waveform_sig_rx =-232;
10858: waveform_sig_rx =-175;
10859: waveform_sig_rx =-450;
10860: waveform_sig_rx =-324;
10861: waveform_sig_rx =-90;
10862: waveform_sig_rx =-399;
10863: waveform_sig_rx =-317;
10864: waveform_sig_rx =-176;
10865: waveform_sig_rx =-182;
10866: waveform_sig_rx =-364;
10867: waveform_sig_rx =-182;
10868: waveform_sig_rx =-114;
10869: waveform_sig_rx =-332;
10870: waveform_sig_rx =-257;
10871: waveform_sig_rx =2;
10872: waveform_sig_rx =-290;
10873: waveform_sig_rx =-318;
10874: waveform_sig_rx =31;
10875: waveform_sig_rx =-238;
10876: waveform_sig_rx =-297;
10877: waveform_sig_rx =-15;
10878: waveform_sig_rx =-127;
10879: waveform_sig_rx =-283;
10880: waveform_sig_rx =-24;
10881: waveform_sig_rx =-276;
10882: waveform_sig_rx =-6;
10883: waveform_sig_rx =-184;
10884: waveform_sig_rx =-52;
10885: waveform_sig_rx =-190;
10886: waveform_sig_rx =-98;
10887: waveform_sig_rx =12;
10888: waveform_sig_rx =-296;
10889: waveform_sig_rx =45;
10890: waveform_sig_rx =-22;
10891: waveform_sig_rx =-290;
10892: waveform_sig_rx =126;
10893: waveform_sig_rx =23;
10894: waveform_sig_rx =-308;
10895: waveform_sig_rx =156;
10896: waveform_sig_rx =26;
10897: waveform_sig_rx =-206;
10898: waveform_sig_rx =100;
10899: waveform_sig_rx =74;
10900: waveform_sig_rx =-145;
10901: waveform_sig_rx =-3;
10902: waveform_sig_rx =172;
10903: waveform_sig_rx =-77;
10904: waveform_sig_rx =5;
10905: waveform_sig_rx =85;
10906: waveform_sig_rx =132;
10907: waveform_sig_rx =-111;
10908: waveform_sig_rx =109;
10909: waveform_sig_rx =224;
10910: waveform_sig_rx =-105;
10911: waveform_sig_rx =92;
10912: waveform_sig_rx =282;
10913: waveform_sig_rx =-75;
10914: waveform_sig_rx =52;
10915: waveform_sig_rx =270;
10916: waveform_sig_rx =39;
10917: waveform_sig_rx =29;
10918: waveform_sig_rx =218;
10919: waveform_sig_rx =189;
10920: waveform_sig_rx =5;
10921: waveform_sig_rx =239;
10922: waveform_sig_rx =64;
10923: waveform_sig_rx =248;
10924: waveform_sig_rx =97;
10925: waveform_sig_rx =293;
10926: waveform_sig_rx =51;
10927: waveform_sig_rx =235;
10928: waveform_sig_rx =325;
10929: waveform_sig_rx =-21;
10930: waveform_sig_rx =362;
10931: waveform_sig_rx =237;
10932: waveform_sig_rx =-24;
10933: waveform_sig_rx =458;
10934: waveform_sig_rx =266;
10935: waveform_sig_rx =-20;
10936: waveform_sig_rx =492;
10937: waveform_sig_rx =249;
10938: waveform_sig_rx =94;
10939: waveform_sig_rx =418;
10940: waveform_sig_rx =318;
10941: waveform_sig_rx =178;
10942: waveform_sig_rx =266;
10943: waveform_sig_rx =449;
10944: waveform_sig_rx =260;
10945: waveform_sig_rx =221;
10946: waveform_sig_rx =418;
10947: waveform_sig_rx =415;
10948: waveform_sig_rx =120;
10949: waveform_sig_rx =469;
10950: waveform_sig_rx =438;
10951: waveform_sig_rx =168;
10952: waveform_sig_rx =414;
10953: waveform_sig_rx =504;
10954: waveform_sig_rx =235;
10955: waveform_sig_rx =334;
10956: waveform_sig_rx =528;
10957: waveform_sig_rx =358;
10958: waveform_sig_rx =290;
10959: waveform_sig_rx =512;
10960: waveform_sig_rx =493;
10961: waveform_sig_rx =297;
10962: waveform_sig_rx =507;
10963: waveform_sig_rx =386;
10964: waveform_sig_rx =511;
10965: waveform_sig_rx =381;
10966: waveform_sig_rx =579;
10967: waveform_sig_rx =284;
10968: waveform_sig_rx =569;
10969: waveform_sig_rx =555;
10970: waveform_sig_rx =214;
10971: waveform_sig_rx =722;
10972: waveform_sig_rx =451;
10973: waveform_sig_rx =288;
10974: waveform_sig_rx =746;
10975: waveform_sig_rx =468;
10976: waveform_sig_rx =319;
10977: waveform_sig_rx =730;
10978: waveform_sig_rx =499;
10979: waveform_sig_rx =410;
10980: waveform_sig_rx =617;
10981: waveform_sig_rx =626;
10982: waveform_sig_rx =439;
10983: waveform_sig_rx =503;
10984: waveform_sig_rx =757;
10985: waveform_sig_rx =478;
10986: waveform_sig_rx =483;
10987: waveform_sig_rx =716;
10988: waveform_sig_rx =632;
10989: waveform_sig_rx =391;
10990: waveform_sig_rx =763;
10991: waveform_sig_rx =654;
10992: waveform_sig_rx =461;
10993: waveform_sig_rx =684;
10994: waveform_sig_rx =740;
10995: waveform_sig_rx =536;
10996: waveform_sig_rx =588;
10997: waveform_sig_rx =775;
10998: waveform_sig_rx =651;
10999: waveform_sig_rx =511;
11000: waveform_sig_rx =791;
11001: waveform_sig_rx =748;
11002: waveform_sig_rx =487;
11003: waveform_sig_rx =825;
11004: waveform_sig_rx =577;
11005: waveform_sig_rx =742;
11006: waveform_sig_rx =686;
11007: waveform_sig_rx =769;
11008: waveform_sig_rx =538;
11009: waveform_sig_rx =863;
11010: waveform_sig_rx =714;
11011: waveform_sig_rx =542;
11012: waveform_sig_rx =964;
11013: waveform_sig_rx =652;
11014: waveform_sig_rx =616;
11015: waveform_sig_rx =947;
11016: waveform_sig_rx =704;
11017: waveform_sig_rx =590;
11018: waveform_sig_rx =935;
11019: waveform_sig_rx =781;
11020: waveform_sig_rx =629;
11021: waveform_sig_rx =842;
11022: waveform_sig_rx =907;
11023: waveform_sig_rx =641;
11024: waveform_sig_rx =758;
11025: waveform_sig_rx =1019;
11026: waveform_sig_rx =670;
11027: waveform_sig_rx =749;
11028: waveform_sig_rx =964;
11029: waveform_sig_rx =814;
11030: waveform_sig_rx =686;
11031: waveform_sig_rx =984;
11032: waveform_sig_rx =858;
11033: waveform_sig_rx =745;
11034: waveform_sig_rx =880;
11035: waveform_sig_rx =994;
11036: waveform_sig_rx =781;
11037: waveform_sig_rx =771;
11038: waveform_sig_rx =1070;
11039: waveform_sig_rx =826;
11040: waveform_sig_rx =721;
11041: waveform_sig_rx =1092;
11042: waveform_sig_rx =878;
11043: waveform_sig_rx =747;
11044: waveform_sig_rx =1069;
11045: waveform_sig_rx =741;
11046: waveform_sig_rx =1001;
11047: waveform_sig_rx =877;
11048: waveform_sig_rx =958;
11049: waveform_sig_rx =814;
11050: waveform_sig_rx =1038;
11051: waveform_sig_rx =919;
11052: waveform_sig_rx =796;
11053: waveform_sig_rx =1120;
11054: waveform_sig_rx =890;
11055: waveform_sig_rx =818;
11056: waveform_sig_rx =1134;
11057: waveform_sig_rx =946;
11058: waveform_sig_rx =800;
11059: waveform_sig_rx =1139;
11060: waveform_sig_rx =991;
11061: waveform_sig_rx =820;
11062: waveform_sig_rx =1063;
11063: waveform_sig_rx =1098;
11064: waveform_sig_rx =762;
11065: waveform_sig_rx =1026;
11066: waveform_sig_rx =1157;
11067: waveform_sig_rx =837;
11068: waveform_sig_rx =995;
11069: waveform_sig_rx =1095;
11070: waveform_sig_rx =1004;
11071: waveform_sig_rx =882;
11072: waveform_sig_rx =1116;
11073: waveform_sig_rx =1075;
11074: waveform_sig_rx =874;
11075: waveform_sig_rx =1026;
11076: waveform_sig_rx =1190;
11077: waveform_sig_rx =865;
11078: waveform_sig_rx =973;
11079: waveform_sig_rx =1234;
11080: waveform_sig_rx =914;
11081: waveform_sig_rx =942;
11082: waveform_sig_rx =1251;
11083: waveform_sig_rx =998;
11084: waveform_sig_rx =961;
11085: waveform_sig_rx =1175;
11086: waveform_sig_rx =922;
11087: waveform_sig_rx =1207;
11088: waveform_sig_rx =976;
11089: waveform_sig_rx =1141;
11090: waveform_sig_rx =936;
11091: waveform_sig_rx =1171;
11092: waveform_sig_rx =1062;
11093: waveform_sig_rx =912;
11094: waveform_sig_rx =1223;
11095: waveform_sig_rx =1050;
11096: waveform_sig_rx =918;
11097: waveform_sig_rx =1283;
11098: waveform_sig_rx =1080;
11099: waveform_sig_rx =847;
11100: waveform_sig_rx =1336;
11101: waveform_sig_rx =1065;
11102: waveform_sig_rx =895;
11103: waveform_sig_rx =1265;
11104: waveform_sig_rx =1125;
11105: waveform_sig_rx =915;
11106: waveform_sig_rx =1197;
11107: waveform_sig_rx =1191;
11108: waveform_sig_rx =1023;
11109: waveform_sig_rx =1072;
11110: waveform_sig_rx =1212;
11111: waveform_sig_rx =1157;
11112: waveform_sig_rx =952;
11113: waveform_sig_rx =1252;
11114: waveform_sig_rx =1148;
11115: waveform_sig_rx =955;
11116: waveform_sig_rx =1165;
11117: waveform_sig_rx =1292;
11118: waveform_sig_rx =967;
11119: waveform_sig_rx =1112;
11120: waveform_sig_rx =1354;
11121: waveform_sig_rx =973;
11122: waveform_sig_rx =1092;
11123: waveform_sig_rx =1298;
11124: waveform_sig_rx =1053;
11125: waveform_sig_rx =1108;
11126: waveform_sig_rx =1157;
11127: waveform_sig_rx =1068;
11128: waveform_sig_rx =1266;
11129: waveform_sig_rx =997;
11130: waveform_sig_rx =1287;
11131: waveform_sig_rx =961;
11132: waveform_sig_rx =1272;
11133: waveform_sig_rx =1178;
11134: waveform_sig_rx =931;
11135: waveform_sig_rx =1369;
11136: waveform_sig_rx =1072;
11137: waveform_sig_rx =963;
11138: waveform_sig_rx =1421;
11139: waveform_sig_rx =1063;
11140: waveform_sig_rx =965;
11141: waveform_sig_rx =1398;
11142: waveform_sig_rx =1058;
11143: waveform_sig_rx =1004;
11144: waveform_sig_rx =1315;
11145: waveform_sig_rx =1144;
11146: waveform_sig_rx =991;
11147: waveform_sig_rx =1204;
11148: waveform_sig_rx =1221;
11149: waveform_sig_rx =1066;
11150: waveform_sig_rx =1062;
11151: waveform_sig_rx =1272;
11152: waveform_sig_rx =1164;
11153: waveform_sig_rx =951;
11154: waveform_sig_rx =1335;
11155: waveform_sig_rx =1174;
11156: waveform_sig_rx =980;
11157: waveform_sig_rx =1244;
11158: waveform_sig_rx =1263;
11159: waveform_sig_rx =976;
11160: waveform_sig_rx =1177;
11161: waveform_sig_rx =1295;
11162: waveform_sig_rx =1026;
11163: waveform_sig_rx =1120;
11164: waveform_sig_rx =1260;
11165: waveform_sig_rx =1121;
11166: waveform_sig_rx =1079;
11167: waveform_sig_rx =1152;
11168: waveform_sig_rx =1134;
11169: waveform_sig_rx =1160;
11170: waveform_sig_rx =1075;
11171: waveform_sig_rx =1284;
11172: waveform_sig_rx =906;
11173: waveform_sig_rx =1372;
11174: waveform_sig_rx =1073;
11175: waveform_sig_rx =980;
11176: waveform_sig_rx =1415;
11177: waveform_sig_rx =968;
11178: waveform_sig_rx =1080;
11179: waveform_sig_rx =1378;
11180: waveform_sig_rx =1021;
11181: waveform_sig_rx =1005;
11182: waveform_sig_rx =1360;
11183: waveform_sig_rx =1058;
11184: waveform_sig_rx =994;
11185: waveform_sig_rx =1295;
11186: waveform_sig_rx =1127;
11187: waveform_sig_rx =1002;
11188: waveform_sig_rx =1181;
11189: waveform_sig_rx =1195;
11190: waveform_sig_rx =1053;
11191: waveform_sig_rx =984;
11192: waveform_sig_rx =1304;
11193: waveform_sig_rx =1089;
11194: waveform_sig_rx =908;
11195: waveform_sig_rx =1367;
11196: waveform_sig_rx =1026;
11197: waveform_sig_rx =979;
11198: waveform_sig_rx =1249;
11199: waveform_sig_rx =1141;
11200: waveform_sig_rx =1008;
11201: waveform_sig_rx =1073;
11202: waveform_sig_rx =1230;
11203: waveform_sig_rx =1034;
11204: waveform_sig_rx =973;
11205: waveform_sig_rx =1289;
11206: waveform_sig_rx =1049;
11207: waveform_sig_rx =990;
11208: waveform_sig_rx =1186;
11209: waveform_sig_rx =993;
11210: waveform_sig_rx =1145;
11211: waveform_sig_rx =1068;
11212: waveform_sig_rx =1147;
11213: waveform_sig_rx =888;
11214: waveform_sig_rx =1295;
11215: waveform_sig_rx =941;
11216: waveform_sig_rx =961;
11217: waveform_sig_rx =1295;
11218: waveform_sig_rx =896;
11219: waveform_sig_rx =1002;
11220: waveform_sig_rx =1273;
11221: waveform_sig_rx =915;
11222: waveform_sig_rx =955;
11223: waveform_sig_rx =1233;
11224: waveform_sig_rx =939;
11225: waveform_sig_rx =957;
11226: waveform_sig_rx =1109;
11227: waveform_sig_rx =1071;
11228: waveform_sig_rx =854;
11229: waveform_sig_rx =1029;
11230: waveform_sig_rx =1169;
11231: waveform_sig_rx =843;
11232: waveform_sig_rx =942;
11233: waveform_sig_rx =1203;
11234: waveform_sig_rx =854;
11235: waveform_sig_rx =926;
11236: waveform_sig_rx =1169;
11237: waveform_sig_rx =918;
11238: waveform_sig_rx =935;
11239: waveform_sig_rx =1004;
11240: waveform_sig_rx =1105;
11241: waveform_sig_rx =845;
11242: waveform_sig_rx =939;
11243: waveform_sig_rx =1177;
11244: waveform_sig_rx =807;
11245: waveform_sig_rx =899;
11246: waveform_sig_rx =1158;
11247: waveform_sig_rx =846;
11248: waveform_sig_rx =914;
11249: waveform_sig_rx =1026;
11250: waveform_sig_rx =859;
11251: waveform_sig_rx =1006;
11252: waveform_sig_rx =878;
11253: waveform_sig_rx =983;
11254: waveform_sig_rx =772;
11255: waveform_sig_rx =1123;
11256: waveform_sig_rx =788;
11257: waveform_sig_rx =854;
11258: waveform_sig_rx =1123;
11259: waveform_sig_rx =735;
11260: waveform_sig_rx =872;
11261: waveform_sig_rx =1041;
11262: waveform_sig_rx =803;
11263: waveform_sig_rx =790;
11264: waveform_sig_rx =1045;
11265: waveform_sig_rx =815;
11266: waveform_sig_rx =750;
11267: waveform_sig_rx =980;
11268: waveform_sig_rx =912;
11269: waveform_sig_rx =612;
11270: waveform_sig_rx =982;
11271: waveform_sig_rx =949;
11272: waveform_sig_rx =650;
11273: waveform_sig_rx =869;
11274: waveform_sig_rx =938;
11275: waveform_sig_rx =748;
11276: waveform_sig_rx =759;
11277: waveform_sig_rx =929;
11278: waveform_sig_rx =818;
11279: waveform_sig_rx =677;
11280: waveform_sig_rx =856;
11281: waveform_sig_rx =929;
11282: waveform_sig_rx =589;
11283: waveform_sig_rx =804;
11284: waveform_sig_rx =948;
11285: waveform_sig_rx =602;
11286: waveform_sig_rx =733;
11287: waveform_sig_rx =949;
11288: waveform_sig_rx =643;
11289: waveform_sig_rx =736;
11290: waveform_sig_rx =790;
11291: waveform_sig_rx =634;
11292: waveform_sig_rx =852;
11293: waveform_sig_rx =658;
11294: waveform_sig_rx =750;
11295: waveform_sig_rx =601;
11296: waveform_sig_rx =896;
11297: waveform_sig_rx =576;
11298: waveform_sig_rx =650;
11299: waveform_sig_rx =837;
11300: waveform_sig_rx =557;
11301: waveform_sig_rx =621;
11302: waveform_sig_rx =852;
11303: waveform_sig_rx =596;
11304: waveform_sig_rx =476;
11305: waveform_sig_rx =925;
11306: waveform_sig_rx =544;
11307: waveform_sig_rx =512;
11308: waveform_sig_rx =844;
11309: waveform_sig_rx =600;
11310: waveform_sig_rx =447;
11311: waveform_sig_rx =759;
11312: waveform_sig_rx =628;
11313: waveform_sig_rx =495;
11314: waveform_sig_rx =583;
11315: waveform_sig_rx =691;
11316: waveform_sig_rx =550;
11317: waveform_sig_rx =465;
11318: waveform_sig_rx =726;
11319: waveform_sig_rx =565;
11320: waveform_sig_rx =402;
11321: waveform_sig_rx =628;
11322: waveform_sig_rx =658;
11323: waveform_sig_rx =320;
11324: waveform_sig_rx =596;
11325: waveform_sig_rx =677;
11326: waveform_sig_rx =317;
11327: waveform_sig_rx =522;
11328: waveform_sig_rx =669;
11329: waveform_sig_rx =374;
11330: waveform_sig_rx =516;
11331: waveform_sig_rx =482;
11332: waveform_sig_rx =434;
11333: waveform_sig_rx =576;
11334: waveform_sig_rx =370;
11335: waveform_sig_rx =568;
11336: waveform_sig_rx =294;
11337: waveform_sig_rx =627;
11338: waveform_sig_rx =362;
11339: waveform_sig_rx =325;
11340: waveform_sig_rx =642;
11341: waveform_sig_rx =296;
11342: waveform_sig_rx =321;
11343: waveform_sig_rx =682;
11344: waveform_sig_rx =243;
11345: waveform_sig_rx =281;
11346: waveform_sig_rx =665;
11347: waveform_sig_rx =197;
11348: waveform_sig_rx =313;
11349: waveform_sig_rx =525;
11350: waveform_sig_rx =318;
11351: waveform_sig_rx =225;
11352: waveform_sig_rx =466;
11353: waveform_sig_rx =368;
11354: waveform_sig_rx =259;
11355: waveform_sig_rx =287;
11356: waveform_sig_rx =446;
11357: waveform_sig_rx =265;
11358: waveform_sig_rx =175;
11359: waveform_sig_rx =474;
11360: waveform_sig_rx =269;
11361: waveform_sig_rx =108;
11362: waveform_sig_rx =438;
11363: waveform_sig_rx =318;
11364: waveform_sig_rx =53;
11365: waveform_sig_rx =353;
11366: waveform_sig_rx =337;
11367: waveform_sig_rx =107;
11368: waveform_sig_rx =225;
11369: waveform_sig_rx =347;
11370: waveform_sig_rx =131;
11371: waveform_sig_rx =194;
11372: waveform_sig_rx =187;
11373: waveform_sig_rx =176;
11374: waveform_sig_rx =225;
11375: waveform_sig_rx =112;
11376: waveform_sig_rx =270;
11377: waveform_sig_rx =-52;
11378: waveform_sig_rx =373;
11379: waveform_sig_rx =31;
11380: waveform_sig_rx =41;
11381: waveform_sig_rx =407;
11382: waveform_sig_rx =-85;
11383: waveform_sig_rx =62;
11384: waveform_sig_rx =381;
11385: waveform_sig_rx =-144;
11386: waveform_sig_rx =69;
11387: waveform_sig_rx =311;
11388: waveform_sig_rx =-115;
11389: waveform_sig_rx =78;
11390: waveform_sig_rx =168;
11391: waveform_sig_rx =61;
11392: waveform_sig_rx =-111;
11393: waveform_sig_rx =128;
11394: waveform_sig_rx =91;
11395: waveform_sig_rx =-99;
11396: waveform_sig_rx =-7;
11397: waveform_sig_rx =174;
11398: waveform_sig_rx =-78;
11399: waveform_sig_rx =-113;
11400: waveform_sig_rx =206;
11401: waveform_sig_rx =-94;
11402: waveform_sig_rx =-172;
11403: waveform_sig_rx =156;
11404: waveform_sig_rx =-35;
11405: waveform_sig_rx =-195;
11406: waveform_sig_rx =30;
11407: waveform_sig_rx =-15;
11408: waveform_sig_rx =-167;
11409: waveform_sig_rx =-144;
11410: waveform_sig_rx =80;
11411: waveform_sig_rx =-187;
11412: waveform_sig_rx =-142;
11413: waveform_sig_rx =-60;
11414: waveform_sig_rx =-167;
11415: waveform_sig_rx =-100;
11416: waveform_sig_rx =-137;
11417: waveform_sig_rx =-109;
11418: waveform_sig_rx =-321;
11419: waveform_sig_rx =102;
11420: waveform_sig_rx =-353;
11421: waveform_sig_rx =-212;
11422: waveform_sig_rx =58;
11423: waveform_sig_rx =-441;
11424: waveform_sig_rx =-146;
11425: waveform_sig_rx =10;
11426: waveform_sig_rx =-438;
11427: waveform_sig_rx =-188;
11428: waveform_sig_rx =-70;
11429: waveform_sig_rx =-378;
11430: waveform_sig_rx =-256;
11431: waveform_sig_rx =-169;
11432: waveform_sig_rx =-202;
11433: waveform_sig_rx =-446;
11434: waveform_sig_rx =-126;
11435: waveform_sig_rx =-202;
11436: waveform_sig_rx =-441;
11437: waveform_sig_rx =-274;
11438: waveform_sig_rx =-152;
11439: waveform_sig_rx =-427;
11440: waveform_sig_rx =-384;
11441: waveform_sig_rx =-129;
11442: waveform_sig_rx =-426;
11443: waveform_sig_rx =-421;
11444: waveform_sig_rx =-174;
11445: waveform_sig_rx =-338;
11446: waveform_sig_rx =-470;
11447: waveform_sig_rx =-317;
11448: waveform_sig_rx =-269;
11449: waveform_sig_rx =-475;
11450: waveform_sig_rx =-479;
11451: waveform_sig_rx =-163;
11452: waveform_sig_rx =-551;
11453: waveform_sig_rx =-434;
11454: waveform_sig_rx =-347;
11455: waveform_sig_rx =-520;
11456: waveform_sig_rx =-371;
11457: waveform_sig_rx =-440;
11458: waveform_sig_rx =-454;
11459: waveform_sig_rx =-540;
11460: waveform_sig_rx =-231;
11461: waveform_sig_rx =-668;
11462: waveform_sig_rx =-430;
11463: waveform_sig_rx =-312;
11464: waveform_sig_rx =-668;
11465: waveform_sig_rx =-436;
11466: waveform_sig_rx =-323;
11467: waveform_sig_rx =-681;
11468: waveform_sig_rx =-521;
11469: waveform_sig_rx =-314;
11470: waveform_sig_rx =-646;
11471: waveform_sig_rx =-552;
11472: waveform_sig_rx =-404;
11473: waveform_sig_rx =-496;
11474: waveform_sig_rx =-751;
11475: waveform_sig_rx =-391;
11476: waveform_sig_rx =-514;
11477: waveform_sig_rx =-712;
11478: waveform_sig_rx =-529;
11479: waveform_sig_rx =-422;
11480: waveform_sig_rx =-712;
11481: waveform_sig_rx =-600;
11482: waveform_sig_rx =-454;
11483: waveform_sig_rx =-703;
11484: waveform_sig_rx =-674;
11485: waveform_sig_rx =-526;
11486: waveform_sig_rx =-537;
11487: waveform_sig_rx =-794;
11488: waveform_sig_rx =-590;
11489: waveform_sig_rx =-486;
11490: waveform_sig_rx =-853;
11491: waveform_sig_rx =-651;
11492: waveform_sig_rx =-454;
11493: waveform_sig_rx =-878;
11494: waveform_sig_rx =-605;
11495: waveform_sig_rx =-715;
11496: waveform_sig_rx =-749;
11497: waveform_sig_rx =-635;
11498: waveform_sig_rx =-772;
11499: waveform_sig_rx =-670;
11500: waveform_sig_rx =-823;
11501: waveform_sig_rx =-542;
11502: waveform_sig_rx =-886;
11503: waveform_sig_rx =-728;
11504: waveform_sig_rx =-592;
11505: waveform_sig_rx =-937;
11506: waveform_sig_rx =-720;
11507: waveform_sig_rx =-585;
11508: waveform_sig_rx =-928;
11509: waveform_sig_rx =-796;
11510: waveform_sig_rx =-568;
11511: waveform_sig_rx =-891;
11512: waveform_sig_rx =-840;
11513: waveform_sig_rx =-633;
11514: waveform_sig_rx =-809;
11515: waveform_sig_rx =-1006;
11516: waveform_sig_rx =-611;
11517: waveform_sig_rx =-837;
11518: waveform_sig_rx =-937;
11519: waveform_sig_rx =-766;
11520: waveform_sig_rx =-731;
11521: waveform_sig_rx =-929;
11522: waveform_sig_rx =-881;
11523: waveform_sig_rx =-712;
11524: waveform_sig_rx =-888;
11525: waveform_sig_rx =-995;
11526: waveform_sig_rx =-723;
11527: waveform_sig_rx =-797;
11528: waveform_sig_rx =-1093;
11529: waveform_sig_rx =-735;
11530: waveform_sig_rx =-802;
11531: waveform_sig_rx =-1090;
11532: waveform_sig_rx =-822;
11533: waveform_sig_rx =-757;
11534: waveform_sig_rx =-1052;
11535: waveform_sig_rx =-827;
11536: waveform_sig_rx =-973;
11537: waveform_sig_rx =-909;
11538: waveform_sig_rx =-898;
11539: waveform_sig_rx =-956;
11540: waveform_sig_rx =-896;
11541: waveform_sig_rx =-1055;
11542: waveform_sig_rx =-729;
11543: waveform_sig_rx =-1114;
11544: waveform_sig_rx =-939;
11545: waveform_sig_rx =-801;
11546: waveform_sig_rx =-1132;
11547: waveform_sig_rx =-946;
11548: waveform_sig_rx =-780;
11549: waveform_sig_rx =-1165;
11550: waveform_sig_rx =-1016;
11551: waveform_sig_rx =-731;
11552: waveform_sig_rx =-1172;
11553: waveform_sig_rx =-1013;
11554: waveform_sig_rx =-800;
11555: waveform_sig_rx =-1105;
11556: waveform_sig_rx =-1127;
11557: waveform_sig_rx =-826;
11558: waveform_sig_rx =-1048;
11559: waveform_sig_rx =-1042;
11560: waveform_sig_rx =-1050;
11561: waveform_sig_rx =-873;
11562: waveform_sig_rx =-1131;
11563: waveform_sig_rx =-1105;
11564: waveform_sig_rx =-831;
11565: waveform_sig_rx =-1141;
11566: waveform_sig_rx =-1147;
11567: waveform_sig_rx =-853;
11568: waveform_sig_rx =-1041;
11569: waveform_sig_rx =-1220;
11570: waveform_sig_rx =-922;
11571: waveform_sig_rx =-988;
11572: waveform_sig_rx =-1216;
11573: waveform_sig_rx =-997;
11574: waveform_sig_rx =-938;
11575: waveform_sig_rx =-1202;
11576: waveform_sig_rx =-989;
11577: waveform_sig_rx =-1138;
11578: waveform_sig_rx =-1029;
11579: waveform_sig_rx =-1088;
11580: waveform_sig_rx =-1069;
11581: waveform_sig_rx =-1048;
11582: waveform_sig_rx =-1224;
11583: waveform_sig_rx =-868;
11584: waveform_sig_rx =-1302;
11585: waveform_sig_rx =-1089;
11586: waveform_sig_rx =-917;
11587: waveform_sig_rx =-1347;
11588: waveform_sig_rx =-1029;
11589: waveform_sig_rx =-904;
11590: waveform_sig_rx =-1345;
11591: waveform_sig_rx =-1061;
11592: waveform_sig_rx =-917;
11593: waveform_sig_rx =-1328;
11594: waveform_sig_rx =-1056;
11595: waveform_sig_rx =-989;
11596: waveform_sig_rx =-1185;
11597: waveform_sig_rx =-1232;
11598: waveform_sig_rx =-994;
11599: waveform_sig_rx =-1111;
11600: waveform_sig_rx =-1227;
11601: waveform_sig_rx =-1132;
11602: waveform_sig_rx =-963;
11603: waveform_sig_rx =-1316;
11604: waveform_sig_rx =-1134;
11605: waveform_sig_rx =-957;
11606: waveform_sig_rx =-1265;
11607: waveform_sig_rx =-1219;
11608: waveform_sig_rx =-982;
11609: waveform_sig_rx =-1189;
11610: waveform_sig_rx =-1289;
11611: waveform_sig_rx =-1011;
11612: waveform_sig_rx =-1121;
11613: waveform_sig_rx =-1272;
11614: waveform_sig_rx =-1114;
11615: waveform_sig_rx =-1010;
11616: waveform_sig_rx =-1236;
11617: waveform_sig_rx =-1128;
11618: waveform_sig_rx =-1165;
11619: waveform_sig_rx =-1105;
11620: waveform_sig_rx =-1205;
11621: waveform_sig_rx =-1062;
11622: waveform_sig_rx =-1196;
11623: waveform_sig_rx =-1232;
11624: waveform_sig_rx =-905;
11625: waveform_sig_rx =-1438;
11626: waveform_sig_rx =-1057;
11627: waveform_sig_rx =-1025;
11628: waveform_sig_rx =-1404;
11629: waveform_sig_rx =-1017;
11630: waveform_sig_rx =-1051;
11631: waveform_sig_rx =-1372;
11632: waveform_sig_rx =-1092;
11633: waveform_sig_rx =-1026;
11634: waveform_sig_rx =-1343;
11635: waveform_sig_rx =-1117;
11636: waveform_sig_rx =-1048;
11637: waveform_sig_rx =-1212;
11638: waveform_sig_rx =-1272;
11639: waveform_sig_rx =-1030;
11640: waveform_sig_rx =-1138;
11641: waveform_sig_rx =-1299;
11642: waveform_sig_rx =-1153;
11643: waveform_sig_rx =-993;
11644: waveform_sig_rx =-1395;
11645: waveform_sig_rx =-1107;
11646: waveform_sig_rx =-1026;
11647: waveform_sig_rx =-1296;
11648: waveform_sig_rx =-1166;
11649: waveform_sig_rx =-1060;
11650: waveform_sig_rx =-1167;
11651: waveform_sig_rx =-1274;
11652: waveform_sig_rx =-1080;
11653: waveform_sig_rx =-1094;
11654: waveform_sig_rx =-1321;
11655: waveform_sig_rx =-1124;
11656: waveform_sig_rx =-986;
11657: waveform_sig_rx =-1332;
11658: waveform_sig_rx =-1085;
11659: waveform_sig_rx =-1160;
11660: waveform_sig_rx =-1161;
11661: waveform_sig_rx =-1144;
11662: waveform_sig_rx =-1083;
11663: waveform_sig_rx =-1238;
11664: waveform_sig_rx =-1148;
11665: waveform_sig_rx =-962;
11666: waveform_sig_rx =-1401;
11667: waveform_sig_rx =-975;
11668: waveform_sig_rx =-1073;
11669: waveform_sig_rx =-1318;
11670: waveform_sig_rx =-1017;
11671: waveform_sig_rx =-1033;
11672: waveform_sig_rx =-1300;
11673: waveform_sig_rx =-1081;
11674: waveform_sig_rx =-967;
11675: waveform_sig_rx =-1295;
11676: waveform_sig_rx =-1102;
11677: waveform_sig_rx =-1007;
11678: waveform_sig_rx =-1171;
11679: waveform_sig_rx =-1261;
11680: waveform_sig_rx =-927;
11681: waveform_sig_rx =-1115;
11682: waveform_sig_rx =-1280;
11683: waveform_sig_rx =-1018;
11684: waveform_sig_rx =-989;
11685: waveform_sig_rx =-1297;
11686: waveform_sig_rx =-994;
11687: waveform_sig_rx =-1051;
11688: waveform_sig_rx =-1164;
11689: waveform_sig_rx =-1142;
11690: waveform_sig_rx =-1012;
11691: waveform_sig_rx =-1028;
11692: waveform_sig_rx =-1301;
11693: waveform_sig_rx =-926;
11694: waveform_sig_rx =-1007;
11695: waveform_sig_rx =-1312;
11696: waveform_sig_rx =-971;
11697: waveform_sig_rx =-972;
11698: waveform_sig_rx =-1256;
11699: waveform_sig_rx =-964;
11700: waveform_sig_rx =-1155;
11701: waveform_sig_rx =-1025;
11702: waveform_sig_rx =-1072;
11703: waveform_sig_rx =-1018;
11704: waveform_sig_rx =-1095;
11705: waveform_sig_rx =-1056;
11706: waveform_sig_rx =-890;
11707: waveform_sig_rx =-1261;
11708: waveform_sig_rx =-904;
11709: waveform_sig_rx =-995;
11710: waveform_sig_rx =-1200;
11711: waveform_sig_rx =-928;
11712: waveform_sig_rx =-933;
11713: waveform_sig_rx =-1165;
11714: waveform_sig_rx =-999;
11715: waveform_sig_rx =-841;
11716: waveform_sig_rx =-1182;
11717: waveform_sig_rx =-1013;
11718: waveform_sig_rx =-829;
11719: waveform_sig_rx =-1127;
11720: waveform_sig_rx =-1116;
11721: waveform_sig_rx =-760;
11722: waveform_sig_rx =-1083;
11723: waveform_sig_rx =-1056;
11724: waveform_sig_rx =-912;
11725: waveform_sig_rx =-904;
11726: waveform_sig_rx =-1087;
11727: waveform_sig_rx =-938;
11728: waveform_sig_rx =-859;
11729: waveform_sig_rx =-1022;
11730: waveform_sig_rx =-1041;
11731: waveform_sig_rx =-776;
11732: waveform_sig_rx =-968;
11733: waveform_sig_rx =-1123;
11734: waveform_sig_rx =-747;
11735: waveform_sig_rx =-927;
11736: waveform_sig_rx =-1093;
11737: waveform_sig_rx =-794;
11738: waveform_sig_rx =-825;
11739: waveform_sig_rx =-1069;
11740: waveform_sig_rx =-779;
11741: waveform_sig_rx =-1020;
11742: waveform_sig_rx =-838;
11743: waveform_sig_rx =-886;
11744: waveform_sig_rx =-856;
11745: waveform_sig_rx =-925;
11746: waveform_sig_rx =-896;
11747: waveform_sig_rx =-739;
11748: waveform_sig_rx =-1053;
11749: waveform_sig_rx =-770;
11750: waveform_sig_rx =-786;
11751: waveform_sig_rx =-1030;
11752: waveform_sig_rx =-765;
11753: waveform_sig_rx =-693;
11754: waveform_sig_rx =-1076;
11755: waveform_sig_rx =-754;
11756: waveform_sig_rx =-659;
11757: waveform_sig_rx =-1060;
11758: waveform_sig_rx =-731;
11759: waveform_sig_rx =-675;
11760: waveform_sig_rx =-961;
11761: waveform_sig_rx =-864;
11762: waveform_sig_rx =-623;
11763: waveform_sig_rx =-884;
11764: waveform_sig_rx =-837;
11765: waveform_sig_rx =-763;
11766: waveform_sig_rx =-676;
11767: waveform_sig_rx =-914;
11768: waveform_sig_rx =-750;
11769: waveform_sig_rx =-608;
11770: waveform_sig_rx =-880;
11771: waveform_sig_rx =-805;
11772: waveform_sig_rx =-539;
11773: waveform_sig_rx =-821;
11774: waveform_sig_rx =-866;
11775: waveform_sig_rx =-555;
11776: waveform_sig_rx =-756;
11777: waveform_sig_rx =-846;
11778: waveform_sig_rx =-611;
11779: waveform_sig_rx =-643;
11780: waveform_sig_rx =-841;
11781: waveform_sig_rx =-585;
11782: waveform_sig_rx =-798;
11783: waveform_sig_rx =-601;
11784: waveform_sig_rx =-737;
11785: waveform_sig_rx =-609;
11786: waveform_sig_rx =-691;
11787: waveform_sig_rx =-707;
11788: waveform_sig_rx =-461;
11789: waveform_sig_rx =-862;
11790: waveform_sig_rx =-531;
11791: waveform_sig_rx =-487;
11792: waveform_sig_rx =-878;
11793: waveform_sig_rx =-445;
11794: waveform_sig_rx =-475;
11795: waveform_sig_rx =-895;
11796: waveform_sig_rx =-425;
11797: waveform_sig_rx =-514;
11798: waveform_sig_rx =-800;
11799: waveform_sig_rx =-469;
11800: waveform_sig_rx =-500;
11801: waveform_sig_rx =-670;
11802: waveform_sig_rx =-637;
11803: waveform_sig_rx =-388;
11804: waveform_sig_rx =-600;
11805: waveform_sig_rx =-621;
11806: waveform_sig_rx =-503;
11807: waveform_sig_rx =-410;
11808: waveform_sig_rx =-695;
11809: waveform_sig_rx =-490;
11810: waveform_sig_rx =-352;
11811: waveform_sig_rx =-679;
11812: waveform_sig_rx =-518;
11813: waveform_sig_rx =-284;
11814: waveform_sig_rx =-608;
11815: waveform_sig_rx =-545;
11816: waveform_sig_rx =-317;
11817: waveform_sig_rx =-503;
11818: waveform_sig_rx =-551;
11819: waveform_sig_rx =-390;
11820: waveform_sig_rx =-327;
11821: waveform_sig_rx =-565;
11822: waveform_sig_rx =-359;
11823: waveform_sig_rx =-470;
11824: waveform_sig_rx =-353;
11825: waveform_sig_rx =-452;
11826: waveform_sig_rx =-294;
11827: waveform_sig_rx =-497;
11828: waveform_sig_rx =-367;
11829: waveform_sig_rx =-212;
11830: waveform_sig_rx =-649;
11831: waveform_sig_rx =-186;
11832: waveform_sig_rx =-296;
11833: waveform_sig_rx =-615;
11834: waveform_sig_rx =-133;
11835: waveform_sig_rx =-301;
11836: waveform_sig_rx =-571;
11837: waveform_sig_rx =-129;
11838: waveform_sig_rx =-283;
11839: waveform_sig_rx =-467;
11840: waveform_sig_rx =-223;
11841: waveform_sig_rx =-234;
11842: waveform_sig_rx =-366;
11843: waveform_sig_rx =-379;
11844: waveform_sig_rx =-105;
11845: waveform_sig_rx =-308;
11846: waveform_sig_rx =-375;
11847: waveform_sig_rx =-174;
11848: waveform_sig_rx =-158;
11849: waveform_sig_rx =-456;
11850: waveform_sig_rx =-159;
11851: waveform_sig_rx =-116;
11852: waveform_sig_rx =-410;
11853: waveform_sig_rx =-210;
11854: waveform_sig_rx =-72;
11855: waveform_sig_rx =-304;
11856: waveform_sig_rx =-270;
11857: waveform_sig_rx =-86;
11858: waveform_sig_rx =-157;
11859: waveform_sig_rx =-303;
11860: waveform_sig_rx =-100;
11861: waveform_sig_rx =-25;
11862: waveform_sig_rx =-343;
11863: waveform_sig_rx =-48;
11864: waveform_sig_rx =-194;
11865: waveform_sig_rx =-102;
11866: waveform_sig_rx =-162;
11867: waveform_sig_rx =-25;
11868: waveform_sig_rx =-245;
11869: waveform_sig_rx =-38;
11870: waveform_sig_rx =14;
11871: waveform_sig_rx =-362;
11872: waveform_sig_rx =140;
11873: waveform_sig_rx =-94;
11874: waveform_sig_rx =-256;
11875: waveform_sig_rx =164;
11876: waveform_sig_rx =-67;
11877: waveform_sig_rx =-227;
11878: waveform_sig_rx =93;
11879: waveform_sig_rx =2;
11880: waveform_sig_rx =-149;
11881: waveform_sig_rx =5;
11882: waveform_sig_rx =120;
11883: waveform_sig_rx =-118;
11884: waveform_sig_rx =-97;
11885: waveform_sig_rx =251;
11886: waveform_sig_rx =-89;
11887: waveform_sig_rx =-61;
11888: waveform_sig_rx =142;
11889: waveform_sig_rx =112;
11890: waveform_sig_rx =-129;
11891: waveform_sig_rx =157;
11892: waveform_sig_rx =144;
11893: waveform_sig_rx =-78;
11894: waveform_sig_rx =102;
11895: waveform_sig_rx =202;
11896: waveform_sig_rx =43;
11897: waveform_sig_rx =5;
11898: waveform_sig_rx =249;
11899: waveform_sig_rx =168;
11900: waveform_sig_rx =-68;
11901: waveform_sig_rx =253;
11902: waveform_sig_rx =246;
11903: waveform_sig_rx =-98;
11904: waveform_sig_rx =328;
11905: waveform_sig_rx =45;
11906: waveform_sig_rx =207;
11907: waveform_sig_rx =192;
11908: waveform_sig_rx =219;
11909: waveform_sig_rx =62;
11910: waveform_sig_rx =283;
11911: waveform_sig_rx =259;
11912: waveform_sig_rx =29;
11913: waveform_sig_rx =391;
11914: waveform_sig_rx =185;
11915: waveform_sig_rx =75;
11916: waveform_sig_rx =391;
11917: waveform_sig_rx =268;
11918: waveform_sig_rx =58;
11919: waveform_sig_rx =388;
11920: waveform_sig_rx =347;
11921: waveform_sig_rx =107;
11922: waveform_sig_rx =333;
11923: waveform_sig_rx =438;
11924: waveform_sig_rx =131;
11925: waveform_sig_rx =253;
11926: waveform_sig_rx =526;
11927: waveform_sig_rx =183;
11928: waveform_sig_rx =265;
11929: waveform_sig_rx =425;
11930: waveform_sig_rx =377;
11931: waveform_sig_rx =205;
11932: waveform_sig_rx =451;
11933: waveform_sig_rx =423;
11934: waveform_sig_rx =261;
11935: waveform_sig_rx =371;
11936: waveform_sig_rx =531;
11937: waveform_sig_rx =330;
11938: waveform_sig_rx =254;
11939: waveform_sig_rx =606;
11940: waveform_sig_rx =387;
11941: waveform_sig_rx =220;
11942: waveform_sig_rx =619;
11943: waveform_sig_rx =432;
11944: waveform_sig_rx =256;
11945: waveform_sig_rx =610;
11946: waveform_sig_rx =253;
11947: waveform_sig_rx =588;
11948: waveform_sig_rx =391;
11949: waveform_sig_rx =489;
11950: waveform_sig_rx =397;
11951: waveform_sig_rx =502;
11952: waveform_sig_rx =568;
11953: waveform_sig_rx =307;
11954: waveform_sig_rx =639;
11955: waveform_sig_rx =519;
11956: waveform_sig_rx =294;
11957: waveform_sig_rx =704;
11958: waveform_sig_rx =557;
11959: waveform_sig_rx =325;
11960: waveform_sig_rx =706;
11961: waveform_sig_rx =615;
11962: waveform_sig_rx =370;
11963: waveform_sig_rx =642;
11964: waveform_sig_rx =709;
11965: waveform_sig_rx =395;
11966: waveform_sig_rx =569;
11967: waveform_sig_rx =787;
11968: waveform_sig_rx =427;
11969: waveform_sig_rx =580;
11970: waveform_sig_rx =660;
11971: waveform_sig_rx =629;
11972: waveform_sig_rx =503;
11973: waveform_sig_rx =653;
11974: waveform_sig_rx =743;
11975: waveform_sig_rx =497;
11976: waveform_sig_rx =595;
11977: waveform_sig_rx =867;
11978: waveform_sig_rx =488;
11979: waveform_sig_rx =569;
11980: waveform_sig_rx =885;
11981: waveform_sig_rx =540;
11982: waveform_sig_rx =569;
11983: waveform_sig_rx =827;
11984: waveform_sig_rx =652;
11985: waveform_sig_rx =587;
11986: waveform_sig_rx =765;
11987: waveform_sig_rx =568;
11988: waveform_sig_rx =819;
11989: waveform_sig_rx =605;
11990: waveform_sig_rx =816;
11991: waveform_sig_rx =602;
11992: waveform_sig_rx =790;
11993: waveform_sig_rx =809;
11994: waveform_sig_rx =524;
11995: waveform_sig_rx =922;
11996: waveform_sig_rx =756;
11997: waveform_sig_rx =577;
11998: waveform_sig_rx =930;
11999: waveform_sig_rx =805;
12000: waveform_sig_rx =537;
12001: waveform_sig_rx =965;
12002: waveform_sig_rx =833;
12003: waveform_sig_rx =536;
12004: waveform_sig_rx =955;
12005: waveform_sig_rx =877;
12006: waveform_sig_rx =604;
12007: waveform_sig_rx =870;
12008: waveform_sig_rx =898;
12009: waveform_sig_rx =741;
12010: waveform_sig_rx =780;
12011: waveform_sig_rx =854;
12012: waveform_sig_rx =936;
12013: waveform_sig_rx =637;
12014: waveform_sig_rx =951;
12015: waveform_sig_rx =977;
12016: waveform_sig_rx =657;
12017: waveform_sig_rx =906;
12018: waveform_sig_rx =1037;
12019: waveform_sig_rx =692;
12020: waveform_sig_rx =841;
12021: waveform_sig_rx =1051;
12022: waveform_sig_rx =780;
12023: waveform_sig_rx =818;
12024: waveform_sig_rx =1012;
12025: waveform_sig_rx =912;
12026: waveform_sig_rx =809;
12027: waveform_sig_rx =964;
12028: waveform_sig_rx =845;
12029: waveform_sig_rx =1014;
12030: waveform_sig_rx =810;
12031: waveform_sig_rx =1055;
12032: waveform_sig_rx =756;
12033: waveform_sig_rx =1024;
12034: waveform_sig_rx =1005;
12035: waveform_sig_rx =720;
12036: waveform_sig_rx =1153;
12037: waveform_sig_rx =925;
12038: waveform_sig_rx =734;
12039: waveform_sig_rx =1209;
12040: waveform_sig_rx =959;
12041: waveform_sig_rx =722;
12042: waveform_sig_rx =1217;
12043: waveform_sig_rx =932;
12044: waveform_sig_rx =804;
12045: waveform_sig_rx =1155;
12046: waveform_sig_rx =979;
12047: waveform_sig_rx =889;
12048: waveform_sig_rx =984;
12049: waveform_sig_rx =1090;
12050: waveform_sig_rx =973;
12051: waveform_sig_rx =877;
12052: waveform_sig_rx =1137;
12053: waveform_sig_rx =1068;
12054: waveform_sig_rx =785;
12055: waveform_sig_rx =1223;
12056: waveform_sig_rx =1039;
12057: waveform_sig_rx =864;
12058: waveform_sig_rx =1108;
12059: waveform_sig_rx =1161;
12060: waveform_sig_rx =899;
12061: waveform_sig_rx =976;
12062: waveform_sig_rx =1211;
12063: waveform_sig_rx =958;
12064: waveform_sig_rx =967;
12065: waveform_sig_rx =1167;
12066: waveform_sig_rx =1060;
12067: waveform_sig_rx =967;
12068: waveform_sig_rx =1110;
12069: waveform_sig_rx =1022;
12070: waveform_sig_rx =1103;
12071: waveform_sig_rx =966;
12072: waveform_sig_rx =1210;
12073: waveform_sig_rx =837;
12074: waveform_sig_rx =1248;
12075: waveform_sig_rx =1084;
12076: waveform_sig_rx =843;
12077: waveform_sig_rx =1355;
12078: waveform_sig_rx =969;
12079: waveform_sig_rx =961;
12080: waveform_sig_rx =1322;
12081: waveform_sig_rx =1008;
12082: waveform_sig_rx =952;
12083: waveform_sig_rx =1280;
12084: waveform_sig_rx =1076;
12085: waveform_sig_rx =980;
12086: waveform_sig_rx =1214;
12087: waveform_sig_rx =1166;
12088: waveform_sig_rx =959;
12089: waveform_sig_rx =1088;
12090: waveform_sig_rx =1261;
12091: waveform_sig_rx =1019;
12092: waveform_sig_rx =1008;
12093: waveform_sig_rx =1277;
12094: waveform_sig_rx =1104;
12095: waveform_sig_rx =919;
12096: waveform_sig_rx =1321;
12097: waveform_sig_rx =1099;
12098: waveform_sig_rx =995;
12099: waveform_sig_rx =1184;
12100: waveform_sig_rx =1212;
12101: waveform_sig_rx =1026;
12102: waveform_sig_rx =1070;
12103: waveform_sig_rx =1276;
12104: waveform_sig_rx =1076;
12105: waveform_sig_rx =1009;
12106: waveform_sig_rx =1291;
12107: waveform_sig_rx =1166;
12108: waveform_sig_rx =979;
12109: waveform_sig_rx =1256;
12110: waveform_sig_rx =1047;
12111: waveform_sig_rx =1190;
12112: waveform_sig_rx =1128;
12113: waveform_sig_rx =1202;
12114: waveform_sig_rx =950;
12115: waveform_sig_rx =1350;
12116: waveform_sig_rx =1050;
12117: waveform_sig_rx =1000;
12118: waveform_sig_rx =1370;
12119: waveform_sig_rx =999;
12120: waveform_sig_rx =1076;
12121: waveform_sig_rx =1330;
12122: waveform_sig_rx =1097;
12123: waveform_sig_rx =1000;
12124: waveform_sig_rx =1317;
12125: waveform_sig_rx =1123;
12126: waveform_sig_rx =1014;
12127: waveform_sig_rx =1255;
12128: waveform_sig_rx =1245;
12129: waveform_sig_rx =981;
12130: waveform_sig_rx =1141;
12131: waveform_sig_rx =1318;
12132: waveform_sig_rx =1001;
12133: waveform_sig_rx =1088;
12134: waveform_sig_rx =1310;
12135: waveform_sig_rx =1098;
12136: waveform_sig_rx =1032;
12137: waveform_sig_rx =1303;
12138: waveform_sig_rx =1132;
12139: waveform_sig_rx =1071;
12140: waveform_sig_rx =1170;
12141: waveform_sig_rx =1288;
12142: waveform_sig_rx =1037;
12143: waveform_sig_rx =1053;
12144: waveform_sig_rx =1361;
12145: waveform_sig_rx =1027;
12146: waveform_sig_rx =1021;
12147: waveform_sig_rx =1351;
12148: waveform_sig_rx =1079;
12149: waveform_sig_rx =1051;
12150: waveform_sig_rx =1269;
12151: waveform_sig_rx =1012;
12152: waveform_sig_rx =1249;
12153: waveform_sig_rx =1084;
12154: waveform_sig_rx =1194;
12155: waveform_sig_rx =1008;
12156: waveform_sig_rx =1299;
12157: waveform_sig_rx =1078;
12158: waveform_sig_rx =1042;
12159: waveform_sig_rx =1301;
12160: waveform_sig_rx =1046;
12161: waveform_sig_rx =1037;
12162: waveform_sig_rx =1310;
12163: waveform_sig_rx =1112;
12164: waveform_sig_rx =958;
12165: waveform_sig_rx =1335;
12166: waveform_sig_rx =1116;
12167: waveform_sig_rx =957;
12168: waveform_sig_rx =1276;
12169: waveform_sig_rx =1215;
12170: waveform_sig_rx =903;
12171: waveform_sig_rx =1197;
12172: waveform_sig_rx =1240;
12173: waveform_sig_rx =960;
12174: waveform_sig_rx =1133;
12175: waveform_sig_rx =1226;
12176: waveform_sig_rx =1094;
12177: waveform_sig_rx =1004;
12178: waveform_sig_rx =1215;
12179: waveform_sig_rx =1145;
12180: waveform_sig_rx =987;
12181: waveform_sig_rx =1127;
12182: waveform_sig_rx =1283;
12183: waveform_sig_rx =908;
12184: waveform_sig_rx =1088;
12185: waveform_sig_rx =1305;
12186: waveform_sig_rx =938;
12187: waveform_sig_rx =1059;
12188: waveform_sig_rx =1256;
12189: waveform_sig_rx =1020;
12190: waveform_sig_rx =1046;
12191: waveform_sig_rx =1147;
12192: waveform_sig_rx =980;
12193: waveform_sig_rx =1196;
12194: waveform_sig_rx =979;
12195: waveform_sig_rx =1161;
12196: waveform_sig_rx =926;
12197: waveform_sig_rx =1210;
12198: waveform_sig_rx =1026;
12199: waveform_sig_rx =903;
12200: waveform_sig_rx =1227;
12201: waveform_sig_rx =991;
12202: waveform_sig_rx =902;
12203: waveform_sig_rx =1247;
12204: waveform_sig_rx =1001;
12205: waveform_sig_rx =820;
12206: waveform_sig_rx =1303;
12207: waveform_sig_rx =957;
12208: waveform_sig_rx =858;
12209: waveform_sig_rx =1228;
12210: waveform_sig_rx =1015;
12211: waveform_sig_rx =846;
12212: waveform_sig_rx =1127;
12213: waveform_sig_rx =1068;
12214: waveform_sig_rx =916;
12215: waveform_sig_rx =960;
12216: waveform_sig_rx =1092;
12217: waveform_sig_rx =1000;
12218: waveform_sig_rx =834;
12219: waveform_sig_rx =1129;
12220: waveform_sig_rx =1006;
12221: waveform_sig_rx =817;
12222: waveform_sig_rx =1067;
12223: waveform_sig_rx =1106;
12224: waveform_sig_rx =780;
12225: waveform_sig_rx =1012;
12226: waveform_sig_rx =1136;
12227: waveform_sig_rx =804;
12228: waveform_sig_rx =931;
12229: waveform_sig_rx =1095;
12230: waveform_sig_rx =889;
12231: waveform_sig_rx =919;
12232: waveform_sig_rx =958;
12233: waveform_sig_rx =875;
12234: waveform_sig_rx =1038;
12235: waveform_sig_rx =823;
12236: waveform_sig_rx =1078;
12237: waveform_sig_rx =731;
12238: waveform_sig_rx =1094;
12239: waveform_sig_rx =896;
12240: waveform_sig_rx =730;
12241: waveform_sig_rx =1161;
12242: waveform_sig_rx =784;
12243: waveform_sig_rx =754;
12244: waveform_sig_rx =1188;
12245: waveform_sig_rx =738;
12246: waveform_sig_rx =754;
12247: waveform_sig_rx =1125;
12248: waveform_sig_rx =732;
12249: waveform_sig_rx =785;
12250: waveform_sig_rx =1020;
12251: waveform_sig_rx =856;
12252: waveform_sig_rx =712;
12253: waveform_sig_rx =921;
12254: waveform_sig_rx =923;
12255: waveform_sig_rx =760;
12256: waveform_sig_rx =776;
12257: waveform_sig_rx =970;
12258: waveform_sig_rx =825;
12259: waveform_sig_rx =658;
12260: waveform_sig_rx =1024;
12261: waveform_sig_rx =803;
12262: waveform_sig_rx =615;
12263: waveform_sig_rx =948;
12264: waveform_sig_rx =833;
12265: waveform_sig_rx =618;
12266: waveform_sig_rx =842;
12267: waveform_sig_rx =864;
12268: waveform_sig_rx =688;
12269: waveform_sig_rx =699;
12270: waveform_sig_rx =897;
12271: waveform_sig_rx =726;
12272: waveform_sig_rx =672;
12273: waveform_sig_rx =796;
12274: waveform_sig_rx =686;
12275: waveform_sig_rx =767;
12276: waveform_sig_rx =680;
12277: waveform_sig_rx =821;
12278: waveform_sig_rx =492;
12279: waveform_sig_rx =946;
12280: waveform_sig_rx =606;
12281: waveform_sig_rx =565;
12282: waveform_sig_rx =968;
12283: waveform_sig_rx =484;
12284: waveform_sig_rx =612;
12285: waveform_sig_rx =922;
12286: waveform_sig_rx =469;
12287: waveform_sig_rx =607;
12288: waveform_sig_rx =847;
12289: waveform_sig_rx =503;
12290: waveform_sig_rx =603;
12291: waveform_sig_rx =716;
12292: waveform_sig_rx =685;
12293: waveform_sig_rx =447;
12294: waveform_sig_rx =675;
12295: waveform_sig_rx =718;
12296: waveform_sig_rx =470;
12297: waveform_sig_rx =567;
12298: waveform_sig_rx =755;
12299: waveform_sig_rx =537;
12300: waveform_sig_rx =454;
12301: waveform_sig_rx =784;
12302: waveform_sig_rx =515;
12303: waveform_sig_rx =421;
12304: waveform_sig_rx =708;
12305: waveform_sig_rx =572;
12306: waveform_sig_rx =448;
12307: waveform_sig_rx =560;
12308: waveform_sig_rx =647;
12309: waveform_sig_rx =464;
12310: waveform_sig_rx =383;
12311: waveform_sig_rx =733;
12312: waveform_sig_rx =430;
12313: waveform_sig_rx =406;
12314: waveform_sig_rx =592;
12315: waveform_sig_rx =369;
12316: waveform_sig_rx =552;
12317: waveform_sig_rx =448;
12318: waveform_sig_rx =514;
12319: waveform_sig_rx =291;
12320: waveform_sig_rx =686;
12321: waveform_sig_rx =300;
12322: waveform_sig_rx =371;
12323: waveform_sig_rx =668;
12324: waveform_sig_rx =212;
12325: waveform_sig_rx =406;
12326: waveform_sig_rx =624;
12327: waveform_sig_rx =239;
12328: waveform_sig_rx =365;
12329: waveform_sig_rx =551;
12330: waveform_sig_rx =281;
12331: waveform_sig_rx =307;
12332: waveform_sig_rx =442;
12333: waveform_sig_rx =451;
12334: waveform_sig_rx =119;
12335: waveform_sig_rx =459;
12336: waveform_sig_rx =443;
12337: waveform_sig_rx =156;
12338: waveform_sig_rx =364;
12339: waveform_sig_rx =449;
12340: waveform_sig_rx =223;
12341: waveform_sig_rx =226;
12342: waveform_sig_rx =457;
12343: waveform_sig_rx =243;
12344: waveform_sig_rx =159;
12345: waveform_sig_rx =371;
12346: waveform_sig_rx =332;
12347: waveform_sig_rx =120;
12348: waveform_sig_rx =272;
12349: waveform_sig_rx =402;
12350: waveform_sig_rx =128;
12351: waveform_sig_rx =134;
12352: waveform_sig_rx =459;
12353: waveform_sig_rx =94;
12354: waveform_sig_rx =180;
12355: waveform_sig_rx =303;
12356: waveform_sig_rx =72;
12357: waveform_sig_rx =294;
12358: waveform_sig_rx =144;
12359: waveform_sig_rx =198;
12360: waveform_sig_rx =47;
12361: waveform_sig_rx =354;
12362: waveform_sig_rx =-7;
12363: waveform_sig_rx =109;
12364: waveform_sig_rx =310;
12365: waveform_sig_rx =-32;
12366: waveform_sig_rx =102;
12367: waveform_sig_rx =293;
12368: waveform_sig_rx =-9;
12369: waveform_sig_rx =-26;
12370: waveform_sig_rx =301;
12371: waveform_sig_rx =-19;
12372: waveform_sig_rx =-22;
12373: waveform_sig_rx =218;
12374: waveform_sig_rx =90;
12375: waveform_sig_rx =-177;
12376: waveform_sig_rx =201;
12377: waveform_sig_rx =76;
12378: waveform_sig_rx =-106;
12379: waveform_sig_rx =48;
12380: waveform_sig_rx =123;
12381: waveform_sig_rx =-64;
12382: waveform_sig_rx =-89;
12383: waveform_sig_rx =124;
12384: waveform_sig_rx =-46;
12385: waveform_sig_rx =-152;
12386: waveform_sig_rx =57;
12387: waveform_sig_rx =45;
12388: waveform_sig_rx =-253;
12389: waveform_sig_rx =-44;
12390: waveform_sig_rx =100;
12391: waveform_sig_rx =-262;
12392: waveform_sig_rx =-102;
12393: waveform_sig_rx =120;
12394: waveform_sig_rx =-262;
12395: waveform_sig_rx =-54;
12396: waveform_sig_rx =-107;
12397: waveform_sig_rx =-185;
12398: waveform_sig_rx =-14;
12399: waveform_sig_rx =-228;
12400: waveform_sig_rx =-69;
12401: waveform_sig_rx =-291;
12402: waveform_sig_rx =19;
12403: waveform_sig_rx =-265;
12404: waveform_sig_rx =-241;
12405: waveform_sig_rx =3;
12406: waveform_sig_rx =-337;
12407: waveform_sig_rx =-242;
12408: waveform_sig_rx =9;
12409: waveform_sig_rx =-364;
12410: waveform_sig_rx =-322;
12411: waveform_sig_rx =19;
12412: waveform_sig_rx =-376;
12413: waveform_sig_rx =-339;
12414: waveform_sig_rx =-89;
12415: waveform_sig_rx =-283;
12416: waveform_sig_rx =-465;
12417: waveform_sig_rx =-104;
12418: waveform_sig_rx =-279;
12419: waveform_sig_rx =-399;
12420: waveform_sig_rx =-285;
12421: waveform_sig_rx =-194;
12422: waveform_sig_rx =-372;
12423: waveform_sig_rx =-411;
12424: waveform_sig_rx =-172;
12425: waveform_sig_rx =-350;
12426: waveform_sig_rx =-490;
12427: waveform_sig_rx =-205;
12428: waveform_sig_rx =-264;
12429: waveform_sig_rx =-577;
12430: waveform_sig_rx =-238;
12431: waveform_sig_rx =-266;
12432: waveform_sig_rx =-534;
12433: waveform_sig_rx =-327;
12434: waveform_sig_rx =-279;
12435: waveform_sig_rx =-503;
12436: waveform_sig_rx =-387;
12437: waveform_sig_rx =-443;
12438: waveform_sig_rx =-396;
12439: waveform_sig_rx =-391;
12440: waveform_sig_rx =-464;
12441: waveform_sig_rx =-342;
12442: waveform_sig_rx =-634;
12443: waveform_sig_rx =-221;
12444: waveform_sig_rx =-605;
12445: waveform_sig_rx =-524;
12446: waveform_sig_rx =-245;
12447: waveform_sig_rx =-669;
12448: waveform_sig_rx =-503;
12449: waveform_sig_rx =-289;
12450: waveform_sig_rx =-674;
12451: waveform_sig_rx =-587;
12452: waveform_sig_rx =-270;
12453: waveform_sig_rx =-689;
12454: waveform_sig_rx =-577;
12455: waveform_sig_rx =-343;
12456: waveform_sig_rx =-611;
12457: waveform_sig_rx =-682;
12458: waveform_sig_rx =-403;
12459: waveform_sig_rx =-570;
12460: waveform_sig_rx =-616;
12461: waveform_sig_rx =-635;
12462: waveform_sig_rx =-413;
12463: waveform_sig_rx =-657;
12464: waveform_sig_rx =-731;
12465: waveform_sig_rx =-349;
12466: waveform_sig_rx =-697;
12467: waveform_sig_rx =-764;
12468: waveform_sig_rx =-417;
12469: waveform_sig_rx =-637;
12470: waveform_sig_rx =-785;
12471: waveform_sig_rx =-534;
12472: waveform_sig_rx =-583;
12473: waveform_sig_rx =-742;
12474: waveform_sig_rx =-677;
12475: waveform_sig_rx =-492;
12476: waveform_sig_rx =-766;
12477: waveform_sig_rx =-699;
12478: waveform_sig_rx =-651;
12479: waveform_sig_rx =-722;
12480: waveform_sig_rx =-690;
12481: waveform_sig_rx =-708;
12482: waveform_sig_rx =-680;
12483: waveform_sig_rx =-872;
12484: waveform_sig_rx =-472;
12485: waveform_sig_rx =-924;
12486: waveform_sig_rx =-753;
12487: waveform_sig_rx =-527;
12488: waveform_sig_rx =-956;
12489: waveform_sig_rx =-749;
12490: waveform_sig_rx =-532;
12491: waveform_sig_rx =-1006;
12492: waveform_sig_rx =-790;
12493: waveform_sig_rx =-556;
12494: waveform_sig_rx =-996;
12495: waveform_sig_rx =-741;
12496: waveform_sig_rx =-691;
12497: waveform_sig_rx =-843;
12498: waveform_sig_rx =-922;
12499: waveform_sig_rx =-750;
12500: waveform_sig_rx =-735;
12501: waveform_sig_rx =-972;
12502: waveform_sig_rx =-851;
12503: waveform_sig_rx =-592;
12504: waveform_sig_rx =-1034;
12505: waveform_sig_rx =-856;
12506: waveform_sig_rx =-629;
12507: waveform_sig_rx =-989;
12508: waveform_sig_rx =-898;
12509: waveform_sig_rx =-736;
12510: waveform_sig_rx =-832;
12511: waveform_sig_rx =-1024;
12512: waveform_sig_rx =-813;
12513: waveform_sig_rx =-779;
12514: waveform_sig_rx =-1024;
12515: waveform_sig_rx =-889;
12516: waveform_sig_rx =-716;
12517: waveform_sig_rx =-1019;
12518: waveform_sig_rx =-908;
12519: waveform_sig_rx =-884;
12520: waveform_sig_rx =-923;
12521: waveform_sig_rx =-924;
12522: waveform_sig_rx =-891;
12523: waveform_sig_rx =-936;
12524: waveform_sig_rx =-1060;
12525: waveform_sig_rx =-695;
12526: waveform_sig_rx =-1170;
12527: waveform_sig_rx =-904;
12528: waveform_sig_rx =-772;
12529: waveform_sig_rx =-1196;
12530: waveform_sig_rx =-870;
12531: waveform_sig_rx =-813;
12532: waveform_sig_rx =-1179;
12533: waveform_sig_rx =-946;
12534: waveform_sig_rx =-829;
12535: waveform_sig_rx =-1131;
12536: waveform_sig_rx =-998;
12537: waveform_sig_rx =-886;
12538: waveform_sig_rx =-987;
12539: waveform_sig_rx =-1181;
12540: waveform_sig_rx =-866;
12541: waveform_sig_rx =-941;
12542: waveform_sig_rx =-1186;
12543: waveform_sig_rx =-968;
12544: waveform_sig_rx =-849;
12545: waveform_sig_rx =-1221;
12546: waveform_sig_rx =-996;
12547: waveform_sig_rx =-895;
12548: waveform_sig_rx =-1121;
12549: waveform_sig_rx =-1081;
12550: waveform_sig_rx =-938;
12551: waveform_sig_rx =-994;
12552: waveform_sig_rx =-1209;
12553: waveform_sig_rx =-956;
12554: waveform_sig_rx =-929;
12555: waveform_sig_rx =-1211;
12556: waveform_sig_rx =-1062;
12557: waveform_sig_rx =-886;
12558: waveform_sig_rx =-1204;
12559: waveform_sig_rx =-1051;
12560: waveform_sig_rx =-1015;
12561: waveform_sig_rx =-1122;
12562: waveform_sig_rx =-1052;
12563: waveform_sig_rx =-1030;
12564: waveform_sig_rx =-1134;
12565: waveform_sig_rx =-1120;
12566: waveform_sig_rx =-893;
12567: waveform_sig_rx =-1334;
12568: waveform_sig_rx =-987;
12569: waveform_sig_rx =-1030;
12570: waveform_sig_rx =-1275;
12571: waveform_sig_rx =-1049;
12572: waveform_sig_rx =-998;
12573: waveform_sig_rx =-1231;
12574: waveform_sig_rx =-1157;
12575: waveform_sig_rx =-907;
12576: waveform_sig_rx =-1275;
12577: waveform_sig_rx =-1148;
12578: waveform_sig_rx =-956;
12579: waveform_sig_rx =-1169;
12580: waveform_sig_rx =-1294;
12581: waveform_sig_rx =-938;
12582: waveform_sig_rx =-1125;
12583: waveform_sig_rx =-1266;
12584: waveform_sig_rx =-1086;
12585: waveform_sig_rx =-989;
12586: waveform_sig_rx =-1279;
12587: waveform_sig_rx =-1099;
12588: waveform_sig_rx =-1025;
12589: waveform_sig_rx =-1212;
12590: waveform_sig_rx =-1201;
12591: waveform_sig_rx =-1046;
12592: waveform_sig_rx =-1067;
12593: waveform_sig_rx =-1346;
12594: waveform_sig_rx =-1036;
12595: waveform_sig_rx =-1008;
12596: waveform_sig_rx =-1358;
12597: waveform_sig_rx =-1076;
12598: waveform_sig_rx =-987;
12599: waveform_sig_rx =-1336;
12600: waveform_sig_rx =-1057;
12601: waveform_sig_rx =-1204;
12602: waveform_sig_rx =-1171;
12603: waveform_sig_rx =-1090;
12604: waveform_sig_rx =-1162;
12605: waveform_sig_rx =-1168;
12606: waveform_sig_rx =-1216;
12607: waveform_sig_rx =-996;
12608: waveform_sig_rx =-1336;
12609: waveform_sig_rx =-1093;
12610: waveform_sig_rx =-1071;
12611: waveform_sig_rx =-1295;
12612: waveform_sig_rx =-1140;
12613: waveform_sig_rx =-999;
12614: waveform_sig_rx =-1328;
12615: waveform_sig_rx =-1188;
12616: waveform_sig_rx =-918;
12617: waveform_sig_rx =-1357;
12618: waveform_sig_rx =-1174;
12619: waveform_sig_rx =-975;
12620: waveform_sig_rx =-1252;
12621: waveform_sig_rx =-1291;
12622: waveform_sig_rx =-955;
12623: waveform_sig_rx =-1209;
12624: waveform_sig_rx =-1254;
12625: waveform_sig_rx =-1123;
12626: waveform_sig_rx =-1067;
12627: waveform_sig_rx =-1276;
12628: waveform_sig_rx =-1166;
12629: waveform_sig_rx =-1025;
12630: waveform_sig_rx =-1216;
12631: waveform_sig_rx =-1265;
12632: waveform_sig_rx =-987;
12633: waveform_sig_rx =-1116;
12634: waveform_sig_rx =-1367;
12635: waveform_sig_rx =-988;
12636: waveform_sig_rx =-1103;
12637: waveform_sig_rx =-1338;
12638: waveform_sig_rx =-1052;
12639: waveform_sig_rx =-1049;
12640: waveform_sig_rx =-1293;
12641: waveform_sig_rx =-1028;
12642: waveform_sig_rx =-1227;
12643: waveform_sig_rx =-1096;
12644: waveform_sig_rx =-1118;
12645: waveform_sig_rx =-1151;
12646: waveform_sig_rx =-1120;
12647: waveform_sig_rx =-1250;
12648: waveform_sig_rx =-949;
12649: waveform_sig_rx =-1317;
12650: waveform_sig_rx =-1125;
12651: waveform_sig_rx =-977;
12652: waveform_sig_rx =-1323;
12653: waveform_sig_rx =-1093;
12654: waveform_sig_rx =-914;
12655: waveform_sig_rx =-1376;
12656: waveform_sig_rx =-1093;
12657: waveform_sig_rx =-909;
12658: waveform_sig_rx =-1348;
12659: waveform_sig_rx =-1066;
12660: waveform_sig_rx =-977;
12661: waveform_sig_rx =-1217;
12662: waveform_sig_rx =-1216;
12663: waveform_sig_rx =-946;
12664: waveform_sig_rx =-1176;
12665: waveform_sig_rx =-1183;
12666: waveform_sig_rx =-1116;
12667: waveform_sig_rx =-986;
12668: waveform_sig_rx =-1223;
12669: waveform_sig_rx =-1135;
12670: waveform_sig_rx =-916;
12671: waveform_sig_rx =-1206;
12672: waveform_sig_rx =-1190;
12673: waveform_sig_rx =-881;
12674: waveform_sig_rx =-1150;
12675: waveform_sig_rx =-1248;
12676: waveform_sig_rx =-895;
12677: waveform_sig_rx =-1086;
12678: waveform_sig_rx =-1198;
12679: waveform_sig_rx =-1009;
12680: waveform_sig_rx =-975;
12681: waveform_sig_rx =-1186;
12682: waveform_sig_rx =-1007;
12683: waveform_sig_rx =-1135;
12684: waveform_sig_rx =-994;
12685: waveform_sig_rx =-1096;
12686: waveform_sig_rx =-1005;
12687: waveform_sig_rx =-1051;
12688: waveform_sig_rx =-1137;
12689: waveform_sig_rx =-805;
12690: waveform_sig_rx =-1271;
12691: waveform_sig_rx =-979;
12692: waveform_sig_rx =-856;
12693: waveform_sig_rx =-1288;
12694: waveform_sig_rx =-903;
12695: waveform_sig_rx =-863;
12696: waveform_sig_rx =-1288;
12697: waveform_sig_rx =-884;
12698: waveform_sig_rx =-883;
12699: waveform_sig_rx =-1209;
12700: waveform_sig_rx =-917;
12701: waveform_sig_rx =-896;
12702: waveform_sig_rx =-1054;
12703: waveform_sig_rx =-1094;
12704: waveform_sig_rx =-828;
12705: waveform_sig_rx =-1000;
12706: waveform_sig_rx =-1061;
12707: waveform_sig_rx =-955;
12708: waveform_sig_rx =-793;
12709: waveform_sig_rx =-1123;
12710: waveform_sig_rx =-954;
12711: waveform_sig_rx =-747;
12712: waveform_sig_rx =-1127;
12713: waveform_sig_rx =-982;
12714: waveform_sig_rx =-736;
12715: waveform_sig_rx =-1036;
12716: waveform_sig_rx =-1028;
12717: waveform_sig_rx =-811;
12718: waveform_sig_rx =-920;
12719: waveform_sig_rx =-1008;
12720: waveform_sig_rx =-912;
12721: waveform_sig_rx =-753;
12722: waveform_sig_rx =-1059;
12723: waveform_sig_rx =-865;
12724: waveform_sig_rx =-915;
12725: waveform_sig_rx =-883;
12726: waveform_sig_rx =-913;
12727: waveform_sig_rx =-794;
12728: waveform_sig_rx =-978;
12729: waveform_sig_rx =-899;
12730: waveform_sig_rx =-660;
12731: waveform_sig_rx =-1150;
12732: waveform_sig_rx =-707;
12733: waveform_sig_rx =-759;
12734: waveform_sig_rx =-1088;
12735: waveform_sig_rx =-674;
12736: waveform_sig_rx =-749;
12737: waveform_sig_rx =-1056;
12738: waveform_sig_rx =-728;
12739: waveform_sig_rx =-725;
12740: waveform_sig_rx =-997;
12741: waveform_sig_rx =-745;
12742: waveform_sig_rx =-721;
12743: waveform_sig_rx =-864;
12744: waveform_sig_rx =-916;
12745: waveform_sig_rx =-627;
12746: waveform_sig_rx =-803;
12747: waveform_sig_rx =-911;
12748: waveform_sig_rx =-737;
12749: waveform_sig_rx =-604;
12750: waveform_sig_rx =-1006;
12751: waveform_sig_rx =-677;
12752: waveform_sig_rx =-619;
12753: waveform_sig_rx =-922;
12754: waveform_sig_rx =-719;
12755: waveform_sig_rx =-660;
12756: waveform_sig_rx =-768;
12757: waveform_sig_rx =-831;
12758: waveform_sig_rx =-645;
12759: waveform_sig_rx =-619;
12760: waveform_sig_rx =-896;
12761: waveform_sig_rx =-638;
12762: waveform_sig_rx =-525;
12763: waveform_sig_rx =-932;
12764: waveform_sig_rx =-554;
12765: waveform_sig_rx =-755;
12766: waveform_sig_rx =-669;
12767: waveform_sig_rx =-654;
12768: waveform_sig_rx =-619;
12769: waveform_sig_rx =-746;
12770: waveform_sig_rx =-646;
12771: waveform_sig_rx =-505;
12772: waveform_sig_rx =-898;
12773: waveform_sig_rx =-474;
12774: waveform_sig_rx =-595;
12775: waveform_sig_rx =-853;
12776: waveform_sig_rx =-458;
12777: waveform_sig_rx =-566;
12778: waveform_sig_rx =-779;
12779: waveform_sig_rx =-494;
12780: waveform_sig_rx =-494;
12781: waveform_sig_rx =-694;
12782: waveform_sig_rx =-590;
12783: waveform_sig_rx =-443;
12784: waveform_sig_rx =-636;
12785: waveform_sig_rx =-708;
12786: waveform_sig_rx =-321;
12787: waveform_sig_rx =-636;
12788: waveform_sig_rx =-652;
12789: waveform_sig_rx =-438;
12790: waveform_sig_rx =-445;
12791: waveform_sig_rx =-677;
12792: waveform_sig_rx =-446;
12793: waveform_sig_rx =-434;
12794: waveform_sig_rx =-595;
12795: waveform_sig_rx =-524;
12796: waveform_sig_rx =-359;
12797: waveform_sig_rx =-486;
12798: waveform_sig_rx =-636;
12799: waveform_sig_rx =-305;
12800: waveform_sig_rx =-412;
12801: waveform_sig_rx =-672;
12802: waveform_sig_rx =-332;
12803: waveform_sig_rx =-342;
12804: waveform_sig_rx =-659;
12805: waveform_sig_rx =-266;
12806: waveform_sig_rx =-553;
12807: waveform_sig_rx =-354;
12808: waveform_sig_rx =-415;
12809: waveform_sig_rx =-392;
12810: waveform_sig_rx =-449;
12811: waveform_sig_rx =-385;
12812: waveform_sig_rx =-248;
12813: waveform_sig_rx =-594;
12814: waveform_sig_rx =-221;
12815: waveform_sig_rx =-317;
12816: waveform_sig_rx =-529;
12817: waveform_sig_rx =-205;
12818: waveform_sig_rx =-267;
12819: waveform_sig_rx =-507;
12820: waveform_sig_rx =-257;
12821: waveform_sig_rx =-212;
12822: waveform_sig_rx =-491;
12823: waveform_sig_rx =-296;
12824: waveform_sig_rx =-108;
12825: waveform_sig_rx =-450;
12826: waveform_sig_rx =-356;
12827: waveform_sig_rx =-56;
12828: waveform_sig_rx =-409;
12829: waveform_sig_rx =-273;
12830: waveform_sig_rx =-226;
12831: waveform_sig_rx =-167;
12832: waveform_sig_rx =-373;
12833: waveform_sig_rx =-236;
12834: waveform_sig_rx =-87;
12835: waveform_sig_rx =-361;
12836: waveform_sig_rx =-273;
12837: waveform_sig_rx =-9;
12838: waveform_sig_rx =-281;
12839: waveform_sig_rx =-321;
12840: waveform_sig_rx =-9;
12841: waveform_sig_rx =-191;
12842: waveform_sig_rx =-336;
12843: waveform_sig_rx =-12;
12844: waveform_sig_rx =-85;
12845: waveform_sig_rx =-334;
12846: waveform_sig_rx =17;
12847: waveform_sig_rx =-283;
12848: waveform_sig_rx =-5;
12849: waveform_sig_rx =-153;
12850: waveform_sig_rx =-84;
12851: waveform_sig_rx =-143;
12852: waveform_sig_rx =-127;
12853: waveform_sig_rx =46;
12854: waveform_sig_rx =-279;
12855: waveform_sig_rx =33;
12856: waveform_sig_rx =28;
12857: waveform_sig_rx =-279;
12858: waveform_sig_rx =76;
12859: waveform_sig_rx =62;
12860: waveform_sig_rx =-319;
12861: waveform_sig_rx =96;
12862: waveform_sig_rx =72;
12863: waveform_sig_rx =-245;
12864: waveform_sig_rx =89;
12865: waveform_sig_rx =99;
12866: waveform_sig_rx =-152;
12867: waveform_sig_rx =-38;
12868: waveform_sig_rx =171;
12869: waveform_sig_rx =-77;
12870: waveform_sig_rx =-21;
12871: waveform_sig_rx =63;
12872: waveform_sig_rx =156;
12873: waveform_sig_rx =-94;
12874: waveform_sig_rx =96;
12875: waveform_sig_rx =208;
12876: waveform_sig_rx =-87;
12877: waveform_sig_rx =50;
12878: waveform_sig_rx =285;
12879: waveform_sig_rx =-28;
12880: waveform_sig_rx =-3;
12881: waveform_sig_rx =321;
12882: waveform_sig_rx =32;
12883: waveform_sig_rx =-10;
12884: waveform_sig_rx =249;
12885: waveform_sig_rx =177;
12886: waveform_sig_rx =33;
12887: waveform_sig_rx =214;
12888: waveform_sig_rx =51;
12889: waveform_sig_rx =258;
12890: waveform_sig_rx =66;
12891: waveform_sig_rx =268;
12892: waveform_sig_rx =84;
12893: waveform_sig_rx =171;
12894: waveform_sig_rx =365;
12895: waveform_sig_rx =-61;
12896: waveform_sig_rx =363;
12897: waveform_sig_rx =292;
12898: waveform_sig_rx =-21;
12899: waveform_sig_rx =433;
12900: waveform_sig_rx =300;
12901: waveform_sig_rx =-20;
12902: waveform_sig_rx =426;
12903: waveform_sig_rx =328;
12904: waveform_sig_rx =65;
12905: waveform_sig_rx =402;
12906: waveform_sig_rx =367;
12907: waveform_sig_rx =167;
12908: waveform_sig_rx =266;
12909: waveform_sig_rx =435;
12910: waveform_sig_rx =269;
12911: waveform_sig_rx =240;
12912: waveform_sig_rx =381;
12913: waveform_sig_rx =479;
12914: waveform_sig_rx =117;
12915: waveform_sig_rx =429;
12916: waveform_sig_rx =477;
12917: waveform_sig_rx =171;
12918: waveform_sig_rx =401;
12919: waveform_sig_rx =519;
12920: waveform_sig_rx =245;
12921: waveform_sig_rx =333;
12922: waveform_sig_rx =517;
12923: waveform_sig_rx =354;
12924: waveform_sig_rx =299;
12925: waveform_sig_rx =476;
12926: waveform_sig_rx =505;
12927: waveform_sig_rx =266;
12928: waveform_sig_rx =482;
12929: waveform_sig_rx =396;
12930: waveform_sig_rx =509;
12931: waveform_sig_rx =400;
12932: waveform_sig_rx =573;
12933: waveform_sig_rx =304;
12934: waveform_sig_rx =549;
12935: waveform_sig_rx =574;
12936: waveform_sig_rx =233;
12937: waveform_sig_rx =687;
12938: waveform_sig_rx =491;
12939: waveform_sig_rx =290;
12940: waveform_sig_rx =714;
12941: waveform_sig_rx =539;
12942: waveform_sig_rx =283;
12943: waveform_sig_rx =713;
12944: waveform_sig_rx =567;
12945: waveform_sig_rx =351;
12946: waveform_sig_rx =674;
12947: waveform_sig_rx =586;
12948: waveform_sig_rx =467;
12949: waveform_sig_rx =500;
12950: waveform_sig_rx =703;
12951: waveform_sig_rx =548;
12952: waveform_sig_rx =440;
12953: waveform_sig_rx =738;
12954: waveform_sig_rx =687;
12955: waveform_sig_rx =351;
12956: waveform_sig_rx =793;
12957: waveform_sig_rx =656;
12958: waveform_sig_rx =475;
12959: waveform_sig_rx =677;
12960: waveform_sig_rx =737;
12961: waveform_sig_rx =584;
12962: waveform_sig_rx =541;
12963: waveform_sig_rx =815;
12964: waveform_sig_rx =647;
12965: waveform_sig_rx =508;
12966: waveform_sig_rx =806;
12967: waveform_sig_rx =730;
12968: waveform_sig_rx =526;
12969: waveform_sig_rx =786;
12970: waveform_sig_rx =617;
12971: waveform_sig_rx =740;
12972: waveform_sig_rx =654;
12973: waveform_sig_rx =803;
12974: waveform_sig_rx =544;
12975: waveform_sig_rx =821;
12976: waveform_sig_rx =772;
12977: waveform_sig_rx =503;
12978: waveform_sig_rx =976;
12979: waveform_sig_rx =695;
12980: waveform_sig_rx =585;
12981: waveform_sig_rx =959;
12982: waveform_sig_rx =741;
12983: waveform_sig_rx =608;
12984: waveform_sig_rx =926;
12985: waveform_sig_rx =809;
12986: waveform_sig_rx =638;
12987: waveform_sig_rx =842;
12988: waveform_sig_rx =906;
12989: waveform_sig_rx =676;
12990: waveform_sig_rx =709;
12991: waveform_sig_rx =1028;
12992: waveform_sig_rx =691;
12993: waveform_sig_rx =714;
12994: waveform_sig_rx =980;
12995: waveform_sig_rx =816;
12996: waveform_sig_rx =680;
12997: waveform_sig_rx =963;
12998: waveform_sig_rx =876;
12999: waveform_sig_rx =750;
13000: waveform_sig_rx =847;
13001: waveform_sig_rx =1007;
13002: waveform_sig_rx =791;
13003: waveform_sig_rx =767;
13004: waveform_sig_rx =1066;
13005: waveform_sig_rx =850;
13006: waveform_sig_rx =758;
13007: waveform_sig_rx =1031;
13008: waveform_sig_rx =945;
13009: waveform_sig_rx =736;
13010: waveform_sig_rx =1023;
13011: waveform_sig_rx =805;
13012: waveform_sig_rx =967;
13013: waveform_sig_rx =906;
13014: waveform_sig_rx =964;
13015: waveform_sig_rx =779;
13016: waveform_sig_rx =1052;
13017: waveform_sig_rx =923;
13018: waveform_sig_rx =776;
13019: waveform_sig_rx =1108;
13020: waveform_sig_rx =888;
13021: waveform_sig_rx =848;
13022: waveform_sig_rx =1088;
13023: waveform_sig_rx =1009;
13024: waveform_sig_rx =758;
13025: waveform_sig_rx =1112;
13026: waveform_sig_rx =1038;
13027: waveform_sig_rx =778;
13028: waveform_sig_rx =1091;
13029: waveform_sig_rx =1081;
13030: waveform_sig_rx =805;
13031: waveform_sig_rx =995;
13032: waveform_sig_rx =1154;
13033: waveform_sig_rx =854;
13034: waveform_sig_rx =951;
13035: waveform_sig_rx =1120;
13036: waveform_sig_rx =1018;
13037: waveform_sig_rx =884;
13038: waveform_sig_rx =1115;
13039: waveform_sig_rx =1075;
13040: waveform_sig_rx =902;
13041: waveform_sig_rx =1004;
13042: waveform_sig_rx =1205;
13043: waveform_sig_rx =916;
13044: waveform_sig_rx =927;
13045: waveform_sig_rx =1248;
13046: waveform_sig_rx =931;
13047: waveform_sig_rx =914;
13048: waveform_sig_rx =1230;
13049: waveform_sig_rx =1028;
13050: waveform_sig_rx =938;
13051: waveform_sig_rx =1184;
13052: waveform_sig_rx =905;
13053: waveform_sig_rx =1187;
13054: waveform_sig_rx =1004;
13055: waveform_sig_rx =1111;
13056: waveform_sig_rx =960;
13057: waveform_sig_rx =1150;
13058: waveform_sig_rx =1088;
13059: waveform_sig_rx =928;
13060: waveform_sig_rx =1204;
13061: waveform_sig_rx =1072;
13062: waveform_sig_rx =905;
13063: waveform_sig_rx =1238;
13064: waveform_sig_rx =1140;
13065: waveform_sig_rx =824;
13066: waveform_sig_rx =1323;
13067: waveform_sig_rx =1093;
13068: waveform_sig_rx =876;
13069: waveform_sig_rx =1261;
13070: waveform_sig_rx =1140;
13071: waveform_sig_rx =932;
13072: waveform_sig_rx =1124;
13073: waveform_sig_rx =1229;
13074: waveform_sig_rx =999;
13075: waveform_sig_rx =1064;
13076: waveform_sig_rx =1215;
13077: waveform_sig_rx =1135;
13078: waveform_sig_rx =952;
13079: waveform_sig_rx =1215;
13080: waveform_sig_rx =1191;
13081: waveform_sig_rx =962;
13082: waveform_sig_rx =1118;
13083: waveform_sig_rx =1310;
13084: waveform_sig_rx =941;
13085: waveform_sig_rx =1075;
13086: waveform_sig_rx =1351;
13087: waveform_sig_rx =976;
13088: waveform_sig_rx =1082;
13089: waveform_sig_rx =1277;
13090: waveform_sig_rx =1104;
13091: waveform_sig_rx =1096;
13092: waveform_sig_rx =1192;
13093: waveform_sig_rx =1047;
13094: waveform_sig_rx =1260;
13095: waveform_sig_rx =1036;
13096: waveform_sig_rx =1254;
13097: waveform_sig_rx =985;
13098: waveform_sig_rx =1222;
13099: waveform_sig_rx =1196;
13100: waveform_sig_rx =951;
13101: waveform_sig_rx =1326;
13102: waveform_sig_rx =1127;
13103: waveform_sig_rx =941;
13104: waveform_sig_rx =1401;
13105: waveform_sig_rx =1142;
13106: waveform_sig_rx =920;
13107: waveform_sig_rx =1421;
13108: waveform_sig_rx =1097;
13109: waveform_sig_rx =984;
13110: waveform_sig_rx =1334;
13111: waveform_sig_rx =1166;
13112: waveform_sig_rx =998;
13113: waveform_sig_rx =1195;
13114: waveform_sig_rx =1242;
13115: waveform_sig_rx =1077;
13116: waveform_sig_rx =1071;
13117: waveform_sig_rx =1223;
13118: waveform_sig_rx =1194;
13119: waveform_sig_rx =968;
13120: waveform_sig_rx =1305;
13121: waveform_sig_rx =1223;
13122: waveform_sig_rx =962;
13123: waveform_sig_rx =1218;
13124: waveform_sig_rx =1300;
13125: waveform_sig_rx =984;
13126: waveform_sig_rx =1149;
13127: waveform_sig_rx =1305;
13128: waveform_sig_rx =1033;
13129: waveform_sig_rx =1082;
13130: waveform_sig_rx =1269;
13131: waveform_sig_rx =1142;
13132: waveform_sig_rx =1050;
13133: waveform_sig_rx =1186;
13134: waveform_sig_rx =1073;
13135: waveform_sig_rx =1217;
13136: waveform_sig_rx =1042;
13137: waveform_sig_rx =1282;
13138: waveform_sig_rx =939;
13139: waveform_sig_rx =1287;
13140: waveform_sig_rx =1174;
13141: waveform_sig_rx =929;
13142: waveform_sig_rx =1389;
13143: waveform_sig_rx =1048;
13144: waveform_sig_rx =993;
13145: waveform_sig_rx =1403;
13146: waveform_sig_rx =1043;
13147: waveform_sig_rx =985;
13148: waveform_sig_rx =1370;
13149: waveform_sig_rx =1056;
13150: waveform_sig_rx =1010;
13151: waveform_sig_rx =1253;
13152: waveform_sig_rx =1172;
13153: waveform_sig_rx =990;
13154: waveform_sig_rx =1154;
13155: waveform_sig_rx =1258;
13156: waveform_sig_rx =1040;
13157: waveform_sig_rx =1048;
13158: waveform_sig_rx =1253;
13159: waveform_sig_rx =1145;
13160: waveform_sig_rx =920;
13161: waveform_sig_rx =1297;
13162: waveform_sig_rx =1137;
13163: waveform_sig_rx =930;
13164: waveform_sig_rx =1225;
13165: waveform_sig_rx =1193;
13166: waveform_sig_rx =984;
13167: waveform_sig_rx =1097;
13168: waveform_sig_rx =1221;
13169: waveform_sig_rx =1053;
13170: waveform_sig_rx =985;
13171: waveform_sig_rx =1262;
13172: waveform_sig_rx =1113;
13173: waveform_sig_rx =950;
13174: waveform_sig_rx =1189;
13175: waveform_sig_rx =1006;
13176: waveform_sig_rx =1150;
13177: waveform_sig_rx =1047;
13178: waveform_sig_rx =1179;
13179: waveform_sig_rx =873;
13180: waveform_sig_rx =1263;
13181: waveform_sig_rx =1014;
13182: waveform_sig_rx =899;
13183: waveform_sig_rx =1310;
13184: waveform_sig_rx =908;
13185: waveform_sig_rx =981;
13186: waveform_sig_rx =1273;
13187: waveform_sig_rx =933;
13188: waveform_sig_rx =928;
13189: waveform_sig_rx =1238;
13190: waveform_sig_rx =991;
13191: waveform_sig_rx =939;
13192: waveform_sig_rx =1134;
13193: waveform_sig_rx =1093;
13194: waveform_sig_rx =861;
13195: waveform_sig_rx =1051;
13196: waveform_sig_rx =1147;
13197: waveform_sig_rx =893;
13198: waveform_sig_rx =958;
13199: waveform_sig_rx =1170;
13200: waveform_sig_rx =973;
13201: waveform_sig_rx =827;
13202: waveform_sig_rx =1202;
13203: waveform_sig_rx =959;
13204: waveform_sig_rx =865;
13205: waveform_sig_rx =1083;
13206: waveform_sig_rx =1035;
13207: waveform_sig_rx =890;
13208: waveform_sig_rx =916;
13209: waveform_sig_rx =1111;
13210: waveform_sig_rx =915;
13211: waveform_sig_rx =794;
13212: waveform_sig_rx =1185;
13213: waveform_sig_rx =897;
13214: waveform_sig_rx =832;
13215: waveform_sig_rx =1096;
13216: waveform_sig_rx =790;
13217: waveform_sig_rx =1048;
13218: waveform_sig_rx =867;
13219: waveform_sig_rx =987;
13220: waveform_sig_rx =771;
13221: waveform_sig_rx =1097;
13222: waveform_sig_rx =856;
13223: waveform_sig_rx =783;
13224: waveform_sig_rx =1122;
13225: waveform_sig_rx =771;
13226: waveform_sig_rx =808;
13227: waveform_sig_rx =1141;
13228: waveform_sig_rx =778;
13229: waveform_sig_rx =782;
13230: waveform_sig_rx =1055;
13231: waveform_sig_rx =817;
13232: waveform_sig_rx =775;
13233: waveform_sig_rx =938;
13234: waveform_sig_rx =966;
13235: waveform_sig_rx =642;
13236: waveform_sig_rx =895;
13237: waveform_sig_rx =982;
13238: waveform_sig_rx =664;
13239: waveform_sig_rx =839;
13240: waveform_sig_rx =969;
13241: waveform_sig_rx =777;
13242: waveform_sig_rx =744;
13243: waveform_sig_rx =960;
13244: waveform_sig_rx =818;
13245: waveform_sig_rx =694;
13246: waveform_sig_rx =851;
13247: waveform_sig_rx =944;
13248: waveform_sig_rx =634;
13249: waveform_sig_rx =748;
13250: waveform_sig_rx =994;
13251: waveform_sig_rx =624;
13252: waveform_sig_rx =690;
13253: waveform_sig_rx =985;
13254: waveform_sig_rx =647;
13255: waveform_sig_rx =725;
13256: waveform_sig_rx =823;
13257: waveform_sig_rx =617;
13258: waveform_sig_rx =860;
13259: waveform_sig_rx =635;
13260: waveform_sig_rx =800;
13261: waveform_sig_rx =550;
13262: waveform_sig_rx =885;
13263: waveform_sig_rx =627;
13264: waveform_sig_rx =590;
13265: waveform_sig_rx =902;
13266: waveform_sig_rx =542;
13267: waveform_sig_rx =619;
13268: waveform_sig_rx =844;
13269: waveform_sig_rx =589;
13270: waveform_sig_rx =544;
13271: waveform_sig_rx =838;
13272: waveform_sig_rx =644;
13273: waveform_sig_rx =480;
13274: waveform_sig_rx =797;
13275: waveform_sig_rx =701;
13276: waveform_sig_rx =384;
13277: waveform_sig_rx =782;
13278: waveform_sig_rx =656;
13279: waveform_sig_rx =499;
13280: waveform_sig_rx =632;
13281: waveform_sig_rx =669;
13282: waveform_sig_rx =611;
13283: waveform_sig_rx =441;
13284: waveform_sig_rx =724;
13285: waveform_sig_rx =610;
13286: waveform_sig_rx =390;
13287: waveform_sig_rx =660;
13288: waveform_sig_rx =667;
13289: waveform_sig_rx =372;
13290: waveform_sig_rx =564;
13291: waveform_sig_rx =688;
13292: waveform_sig_rx =407;
13293: waveform_sig_rx =458;
13294: waveform_sig_rx =705;
13295: waveform_sig_rx =408;
13296: waveform_sig_rx =464;
13297: waveform_sig_rx =555;
13298: waveform_sig_rx =391;
13299: waveform_sig_rx =593;
13300: waveform_sig_rx =384;
13301: waveform_sig_rx =569;
13302: waveform_sig_rx =303;
13303: waveform_sig_rx =621;
13304: waveform_sig_rx =389;
13305: waveform_sig_rx =326;
13306: waveform_sig_rx =611;
13307: waveform_sig_rx =317;
13308: waveform_sig_rx =295;
13309: waveform_sig_rx =652;
13310: waveform_sig_rx =303;
13311: waveform_sig_rx =226;
13312: waveform_sig_rx =656;
13313: waveform_sig_rx =259;
13314: waveform_sig_rx =265;
13315: waveform_sig_rx =564;
13316: waveform_sig_rx =347;
13317: waveform_sig_rx =219;
13318: waveform_sig_rx =465;
13319: waveform_sig_rx =376;
13320: waveform_sig_rx =291;
13321: waveform_sig_rx =271;
13322: waveform_sig_rx =481;
13323: waveform_sig_rx =293;
13324: waveform_sig_rx =146;
13325: waveform_sig_rx =517;
13326: waveform_sig_rx =246;
13327: waveform_sig_rx =132;
13328: waveform_sig_rx =386;
13329: waveform_sig_rx =340;
13330: waveform_sig_rx =83;
13331: waveform_sig_rx =278;
13332: waveform_sig_rx =393;
13333: waveform_sig_rx =83;
13334: waveform_sig_rx =199;
13335: waveform_sig_rx =373;
13336: waveform_sig_rx =123;
13337: waveform_sig_rx =234;
13338: waveform_sig_rx =210;
13339: waveform_sig_rx =167;
13340: waveform_sig_rx =278;
13341: waveform_sig_rx =100;
13342: waveform_sig_rx =307;
13343: waveform_sig_rx =-40;
13344: waveform_sig_rx =361;
13345: waveform_sig_rx =78;
13346: waveform_sig_rx =3;
13347: waveform_sig_rx =377;
13348: waveform_sig_rx =-49;
13349: waveform_sig_rx =41;
13350: waveform_sig_rx =377;
13351: waveform_sig_rx =-93;
13352: waveform_sig_rx =25;
13353: waveform_sig_rx =302;
13354: waveform_sig_rx =-64;
13355: waveform_sig_rx =16;
13356: waveform_sig_rx =182;
13357: waveform_sig_rx =52;
13358: waveform_sig_rx =-108;
13359: waveform_sig_rx =132;
13360: waveform_sig_rx =112;
13361: waveform_sig_rx =-84;
13362: waveform_sig_rx =-27;
13363: waveform_sig_rx =178;
13364: waveform_sig_rx =-58;
13365: waveform_sig_rx =-124;
13366: waveform_sig_rx =194;
13367: waveform_sig_rx =-62;
13368: waveform_sig_rx =-167;
13369: waveform_sig_rx =114;
13370: waveform_sig_rx =13;
13371: waveform_sig_rx =-211;
13372: waveform_sig_rx =20;
13373: waveform_sig_rx =37;
13374: waveform_sig_rx =-188;
13375: waveform_sig_rx =-119;
13376: waveform_sig_rx =84;
13377: waveform_sig_rx =-160;
13378: waveform_sig_rx =-159;
13379: waveform_sig_rx =-56;
13380: waveform_sig_rx =-153;
13381: waveform_sig_rx =-96;
13382: waveform_sig_rx =-142;
13383: waveform_sig_rx =-76;
13384: waveform_sig_rx =-334;
13385: waveform_sig_rx =94;
13386: waveform_sig_rx =-319;
13387: waveform_sig_rx =-247;
13388: waveform_sig_rx =63;
13389: waveform_sig_rx =-386;
13390: waveform_sig_rx =-196;
13391: waveform_sig_rx =26;
13392: waveform_sig_rx =-375;
13393: waveform_sig_rx =-269;
13394: waveform_sig_rx =-19;
13395: waveform_sig_rx =-376;
13396: waveform_sig_rx =-281;
13397: waveform_sig_rx =-148;
13398: waveform_sig_rx =-243;
13399: waveform_sig_rx =-418;
13400: waveform_sig_rx =-192;
13401: waveform_sig_rx =-184;
13402: waveform_sig_rx =-404;
13403: waveform_sig_rx =-332;
13404: waveform_sig_rx =-104;
13405: waveform_sig_rx =-426;
13406: waveform_sig_rx =-393;
13407: waveform_sig_rx =-127;
13408: waveform_sig_rx =-415;
13409: waveform_sig_rx =-417;
13410: waveform_sig_rx =-247;
13411: waveform_sig_rx =-301;
13412: waveform_sig_rx =-487;
13413: waveform_sig_rx =-363;
13414: waveform_sig_rx =-235;
13415: waveform_sig_rx =-494;
13416: waveform_sig_rx =-462;
13417: waveform_sig_rx =-181;
13418: waveform_sig_rx =-504;
13419: waveform_sig_rx =-434;
13420: waveform_sig_rx =-353;
13421: waveform_sig_rx =-498;
13422: waveform_sig_rx =-364;
13423: waveform_sig_rx =-446;
13424: waveform_sig_rx =-414;
13425: waveform_sig_rx =-576;
13426: waveform_sig_rx =-214;
13427: waveform_sig_rx =-640;
13428: waveform_sig_rx =-468;
13429: waveform_sig_rx =-287;
13430: waveform_sig_rx =-658;
13431: waveform_sig_rx =-489;
13432: waveform_sig_rx =-314;
13433: waveform_sig_rx =-647;
13434: waveform_sig_rx =-572;
13435: waveform_sig_rx =-320;
13436: waveform_sig_rx =-652;
13437: waveform_sig_rx =-576;
13438: waveform_sig_rx =-446;
13439: waveform_sig_rx =-513;
13440: waveform_sig_rx =-738;
13441: waveform_sig_rx =-427;
13442: waveform_sig_rx =-465;
13443: waveform_sig_rx =-739;
13444: waveform_sig_rx =-540;
13445: waveform_sig_rx =-427;
13446: waveform_sig_rx =-719;
13447: waveform_sig_rx =-602;
13448: waveform_sig_rx =-475;
13449: waveform_sig_rx =-649;
13450: waveform_sig_rx =-712;
13451: waveform_sig_rx =-552;
13452: waveform_sig_rx =-515;
13453: waveform_sig_rx =-828;
13454: waveform_sig_rx =-584;
13455: waveform_sig_rx =-498;
13456: waveform_sig_rx =-825;
13457: waveform_sig_rx =-675;
13458: waveform_sig_rx =-490;
13459: waveform_sig_rx =-800;
13460: waveform_sig_rx =-691;
13461: waveform_sig_rx =-663;
13462: waveform_sig_rx =-756;
13463: waveform_sig_rx =-625;
13464: waveform_sig_rx =-726;
13465: waveform_sig_rx =-699;
13466: waveform_sig_rx =-819;
13467: waveform_sig_rx =-536;
13468: waveform_sig_rx =-914;
13469: waveform_sig_rx =-729;
13470: waveform_sig_rx =-605;
13471: waveform_sig_rx =-893;
13472: waveform_sig_rx =-777;
13473: waveform_sig_rx =-582;
13474: waveform_sig_rx =-875;
13475: waveform_sig_rx =-884;
13476: waveform_sig_rx =-532;
13477: waveform_sig_rx =-914;
13478: waveform_sig_rx =-860;
13479: waveform_sig_rx =-626;
13480: waveform_sig_rx =-806;
13481: waveform_sig_rx =-975;
13482: waveform_sig_rx =-647;
13483: waveform_sig_rx =-776;
13484: waveform_sig_rx =-947;
13485: waveform_sig_rx =-790;
13486: waveform_sig_rx =-698;
13487: waveform_sig_rx =-930;
13488: waveform_sig_rx =-865;
13489: waveform_sig_rx =-720;
13490: waveform_sig_rx =-870;
13491: waveform_sig_rx =-963;
13492: waveform_sig_rx =-744;
13493: waveform_sig_rx =-758;
13494: waveform_sig_rx =-1085;
13495: waveform_sig_rx =-754;
13496: waveform_sig_rx =-739;
13497: waveform_sig_rx =-1072;
13498: waveform_sig_rx =-846;
13499: waveform_sig_rx =-732;
13500: waveform_sig_rx =-1041;
13501: waveform_sig_rx =-846;
13502: waveform_sig_rx =-929;
13503: waveform_sig_rx =-935;
13504: waveform_sig_rx =-850;
13505: waveform_sig_rx =-983;
13506: waveform_sig_rx =-877;
13507: waveform_sig_rx =-1044;
13508: waveform_sig_rx =-749;
13509: waveform_sig_rx =-1067;
13510: waveform_sig_rx =-975;
13511: waveform_sig_rx =-787;
13512: waveform_sig_rx =-1100;
13513: waveform_sig_rx =-1009;
13514: waveform_sig_rx =-729;
13515: waveform_sig_rx =-1138;
13516: waveform_sig_rx =-1045;
13517: waveform_sig_rx =-710;
13518: waveform_sig_rx =-1182;
13519: waveform_sig_rx =-1012;
13520: waveform_sig_rx =-825;
13521: waveform_sig_rx =-1043;
13522: waveform_sig_rx =-1153;
13523: waveform_sig_rx =-851;
13524: waveform_sig_rx =-988;
13525: waveform_sig_rx =-1105;
13526: waveform_sig_rx =-1007;
13527: waveform_sig_rx =-885;
13528: waveform_sig_rx =-1128;
13529: waveform_sig_rx =-1092;
13530: waveform_sig_rx =-875;
13531: waveform_sig_rx =-1072;
13532: waveform_sig_rx =-1188;
13533: waveform_sig_rx =-879;
13534: waveform_sig_rx =-977;
13535: waveform_sig_rx =-1265;
13536: waveform_sig_rx =-899;
13537: waveform_sig_rx =-987;
13538: waveform_sig_rx =-1206;
13539: waveform_sig_rx =-1005;
13540: waveform_sig_rx =-938;
13541: waveform_sig_rx =-1146;
13542: waveform_sig_rx =-1018;
13543: waveform_sig_rx =-1088;
13544: waveform_sig_rx =-1044;
13545: waveform_sig_rx =-1057;
13546: waveform_sig_rx =-1093;
13547: waveform_sig_rx =-1013;
13548: waveform_sig_rx =-1232;
13549: waveform_sig_rx =-858;
13550: waveform_sig_rx =-1246;
13551: waveform_sig_rx =-1116;
13552: waveform_sig_rx =-878;
13553: waveform_sig_rx =-1308;
13554: waveform_sig_rx =-1107;
13555: waveform_sig_rx =-876;
13556: waveform_sig_rx =-1336;
13557: waveform_sig_rx =-1112;
13558: waveform_sig_rx =-896;
13559: waveform_sig_rx =-1325;
13560: waveform_sig_rx =-1109;
13561: waveform_sig_rx =-994;
13562: waveform_sig_rx =-1173;
13563: waveform_sig_rx =-1253;
13564: waveform_sig_rx =-989;
13565: waveform_sig_rx =-1106;
13566: waveform_sig_rx =-1218;
13567: waveform_sig_rx =-1146;
13568: waveform_sig_rx =-963;
13569: waveform_sig_rx =-1248;
13570: waveform_sig_rx =-1207;
13571: waveform_sig_rx =-927;
13572: waveform_sig_rx =-1232;
13573: waveform_sig_rx =-1243;
13574: waveform_sig_rx =-952;
13575: waveform_sig_rx =-1161;
13576: waveform_sig_rx =-1287;
13577: waveform_sig_rx =-1018;
13578: waveform_sig_rx =-1098;
13579: waveform_sig_rx =-1248;
13580: waveform_sig_rx =-1142;
13581: waveform_sig_rx =-995;
13582: waveform_sig_rx =-1267;
13583: waveform_sig_rx =-1121;
13584: waveform_sig_rx =-1157;
13585: waveform_sig_rx =-1158;
13586: waveform_sig_rx =-1156;
13587: waveform_sig_rx =-1132;
13588: waveform_sig_rx =-1149;
13589: waveform_sig_rx =-1281;
13590: waveform_sig_rx =-901;
13591: waveform_sig_rx =-1367;
13592: waveform_sig_rx =-1149;
13593: waveform_sig_rx =-958;
13594: waveform_sig_rx =-1424;
13595: waveform_sig_rx =-1082;
13596: waveform_sig_rx =-981;
13597: waveform_sig_rx =-1395;
13598: waveform_sig_rx =-1096;
13599: waveform_sig_rx =-1004;
13600: waveform_sig_rx =-1338;
13601: waveform_sig_rx =-1133;
13602: waveform_sig_rx =-1050;
13603: waveform_sig_rx =-1167;
13604: waveform_sig_rx =-1300;
13605: waveform_sig_rx =-1010;
13606: waveform_sig_rx =-1126;
13607: waveform_sig_rx =-1277;
13608: waveform_sig_rx =-1149;
13609: waveform_sig_rx =-986;
13610: waveform_sig_rx =-1319;
13611: waveform_sig_rx =-1166;
13612: waveform_sig_rx =-981;
13613: waveform_sig_rx =-1287;
13614: waveform_sig_rx =-1203;
13615: waveform_sig_rx =-1018;
13616: waveform_sig_rx =-1165;
13617: waveform_sig_rx =-1286;
13618: waveform_sig_rx =-1061;
13619: waveform_sig_rx =-1083;
13620: waveform_sig_rx =-1283;
13621: waveform_sig_rx =-1155;
13622: waveform_sig_rx =-966;
13623: waveform_sig_rx =-1303;
13624: waveform_sig_rx =-1140;
13625: waveform_sig_rx =-1159;
13626: waveform_sig_rx =-1155;
13627: waveform_sig_rx =-1139;
13628: waveform_sig_rx =-1116;
13629: waveform_sig_rx =-1175;
13630: waveform_sig_rx =-1218;
13631: waveform_sig_rx =-908;
13632: waveform_sig_rx =-1380;
13633: waveform_sig_rx =-1042;
13634: waveform_sig_rx =-1008;
13635: waveform_sig_rx =-1360;
13636: waveform_sig_rx =-1007;
13637: waveform_sig_rx =-1008;
13638: waveform_sig_rx =-1300;
13639: waveform_sig_rx =-1093;
13640: waveform_sig_rx =-973;
13641: waveform_sig_rx =-1268;
13642: waveform_sig_rx =-1127;
13643: waveform_sig_rx =-975;
13644: waveform_sig_rx =-1149;
13645: waveform_sig_rx =-1276;
13646: waveform_sig_rx =-925;
13647: waveform_sig_rx =-1113;
13648: waveform_sig_rx =-1232;
13649: waveform_sig_rx =-1071;
13650: waveform_sig_rx =-964;
13651: waveform_sig_rx =-1284;
13652: waveform_sig_rx =-1087;
13653: waveform_sig_rx =-942;
13654: waveform_sig_rx =-1205;
13655: waveform_sig_rx =-1117;
13656: waveform_sig_rx =-1003;
13657: waveform_sig_rx =-1067;
13658: waveform_sig_rx =-1219;
13659: waveform_sig_rx =-1012;
13660: waveform_sig_rx =-954;
13661: waveform_sig_rx =-1276;
13662: waveform_sig_rx =-1026;
13663: waveform_sig_rx =-891;
13664: waveform_sig_rx =-1280;
13665: waveform_sig_rx =-930;
13666: waveform_sig_rx =-1132;
13667: waveform_sig_rx =-1044;
13668: waveform_sig_rx =-1007;
13669: waveform_sig_rx =-1062;
13670: waveform_sig_rx =-1056;
13671: waveform_sig_rx =-1091;
13672: waveform_sig_rx =-856;
13673: waveform_sig_rx =-1237;
13674: waveform_sig_rx =-949;
13675: waveform_sig_rx =-924;
13676: waveform_sig_rx =-1226;
13677: waveform_sig_rx =-932;
13678: waveform_sig_rx =-901;
13679: waveform_sig_rx =-1208;
13680: waveform_sig_rx =-971;
13681: waveform_sig_rx =-850;
13682: waveform_sig_rx =-1161;
13683: waveform_sig_rx =-1030;
13684: waveform_sig_rx =-849;
13685: waveform_sig_rx =-1040;
13686: waveform_sig_rx =-1142;
13687: waveform_sig_rx =-769;
13688: waveform_sig_rx =-1024;
13689: waveform_sig_rx =-1082;
13690: waveform_sig_rx =-912;
13691: waveform_sig_rx =-860;
13692: waveform_sig_rx =-1097;
13693: waveform_sig_rx =-938;
13694: waveform_sig_rx =-838;
13695: waveform_sig_rx =-1009;
13696: waveform_sig_rx =-1004;
13697: waveform_sig_rx =-797;
13698: waveform_sig_rx =-897;
13699: waveform_sig_rx =-1134;
13700: waveform_sig_rx =-788;
13701: waveform_sig_rx =-848;
13702: waveform_sig_rx =-1137;
13703: waveform_sig_rx =-796;
13704: waveform_sig_rx =-818;
13705: waveform_sig_rx =-1095;
13706: waveform_sig_rx =-761;
13707: waveform_sig_rx =-1034;
13708: waveform_sig_rx =-822;
13709: waveform_sig_rx =-913;
13710: waveform_sig_rx =-873;
13711: waveform_sig_rx =-876;
13712: waveform_sig_rx =-967;
13713: waveform_sig_rx =-678;
13714: waveform_sig_rx =-1075;
13715: waveform_sig_rx =-779;
13716: waveform_sig_rx =-743;
13717: waveform_sig_rx =-1056;
13718: waveform_sig_rx =-725;
13719: waveform_sig_rx =-727;
13720: waveform_sig_rx =-1018;
13721: waveform_sig_rx =-798;
13722: waveform_sig_rx =-646;
13723: waveform_sig_rx =-1000;
13724: waveform_sig_rx =-834;
13725: waveform_sig_rx =-601;
13726: waveform_sig_rx =-936;
13727: waveform_sig_rx =-918;
13728: waveform_sig_rx =-573;
13729: waveform_sig_rx =-917;
13730: waveform_sig_rx =-796;
13731: waveform_sig_rx =-770;
13732: waveform_sig_rx =-669;
13733: waveform_sig_rx =-886;
13734: waveform_sig_rx =-817;
13735: waveform_sig_rx =-557;
13736: waveform_sig_rx =-869;
13737: waveform_sig_rx =-823;
13738: waveform_sig_rx =-523;
13739: waveform_sig_rx =-798;
13740: waveform_sig_rx =-854;
13741: waveform_sig_rx =-558;
13742: waveform_sig_rx =-698;
13743: waveform_sig_rx =-876;
13744: waveform_sig_rx =-626;
13745: waveform_sig_rx =-605;
13746: waveform_sig_rx =-850;
13747: waveform_sig_rx =-586;
13748: waveform_sig_rx =-788;
13749: waveform_sig_rx =-608;
13750: waveform_sig_rx =-694;
13751: waveform_sig_rx =-636;
13752: waveform_sig_rx =-673;
13753: waveform_sig_rx =-736;
13754: waveform_sig_rx =-467;
13755: waveform_sig_rx =-851;
13756: waveform_sig_rx =-569;
13757: waveform_sig_rx =-498;
13758: waveform_sig_rx =-844;
13759: waveform_sig_rx =-537;
13760: waveform_sig_rx =-451;
13761: waveform_sig_rx =-866;
13762: waveform_sig_rx =-515;
13763: waveform_sig_rx =-419;
13764: waveform_sig_rx =-832;
13765: waveform_sig_rx =-504;
13766: waveform_sig_rx =-462;
13767: waveform_sig_rx =-679;
13768: waveform_sig_rx =-610;
13769: waveform_sig_rx =-422;
13770: waveform_sig_rx =-568;
13771: waveform_sig_rx =-608;
13772: waveform_sig_rx =-547;
13773: waveform_sig_rx =-339;
13774: waveform_sig_rx =-701;
13775: waveform_sig_rx =-485;
13776: waveform_sig_rx =-331;
13777: waveform_sig_rx =-680;
13778: waveform_sig_rx =-518;
13779: waveform_sig_rx =-325;
13780: waveform_sig_rx =-539;
13781: waveform_sig_rx =-591;
13782: waveform_sig_rx =-326;
13783: waveform_sig_rx =-441;
13784: waveform_sig_rx =-601;
13785: waveform_sig_rx =-343;
13786: waveform_sig_rx =-325;
13787: waveform_sig_rx =-571;
13788: waveform_sig_rx =-335;
13789: waveform_sig_rx =-516;
13790: waveform_sig_rx =-314;
13791: waveform_sig_rx =-466;
13792: waveform_sig_rx =-320;
13793: waveform_sig_rx =-438;
13794: waveform_sig_rx =-461;
13795: waveform_sig_rx =-143;
13796: waveform_sig_rx =-633;
13797: waveform_sig_rx =-260;
13798: waveform_sig_rx =-228;
13799: waveform_sig_rx =-622;
13800: waveform_sig_rx =-177;
13801: waveform_sig_rx =-236;
13802: waveform_sig_rx =-587;
13803: waveform_sig_rx =-174;
13804: waveform_sig_rx =-237;
13805: waveform_sig_rx =-493;
13806: waveform_sig_rx =-234;
13807: waveform_sig_rx =-234;
13808: waveform_sig_rx =-347;
13809: waveform_sig_rx =-406;
13810: waveform_sig_rx =-120;
13811: waveform_sig_rx =-292;
13812: waveform_sig_rx =-388;
13813: waveform_sig_rx =-187;
13814: waveform_sig_rx =-132;
13815: waveform_sig_rx =-437;
13816: waveform_sig_rx =-146;
13817: waveform_sig_rx =-99;
13818: waveform_sig_rx =-349;
13819: waveform_sig_rx =-221;
13820: waveform_sig_rx =-35;
13821: waveform_sig_rx =-255;
13822: waveform_sig_rx =-295;
13823: waveform_sig_rx =-29;
13824: waveform_sig_rx =-184;
13825: waveform_sig_rx =-272;
13826: waveform_sig_rx =-110;
13827: waveform_sig_rx =-45;
13828: waveform_sig_rx =-277;
13829: waveform_sig_rx =-89;
13830: waveform_sig_rx =-163;
13831: waveform_sig_rx =-80;
13832: waveform_sig_rx =-170;
13833: waveform_sig_rx =-12;
13834: waveform_sig_rx =-241;
13835: waveform_sig_rx =-77;
13836: waveform_sig_rx =68;
13837: waveform_sig_rx =-363;
13838: waveform_sig_rx =117;
13839: waveform_sig_rx =-62;
13840: waveform_sig_rx =-265;
13841: waveform_sig_rx =115;
13842: waveform_sig_rx =2;
13843: waveform_sig_rx =-235;
13844: waveform_sig_rx =60;
13845: waveform_sig_rx =79;
13846: waveform_sig_rx =-206;
13847: waveform_sig_rx =24;
13848: waveform_sig_rx =89;
13849: waveform_sig_rx =-83;
13850: waveform_sig_rx =-97;
13851: waveform_sig_rx =184;
13852: waveform_sig_rx =-23;
13853: waveform_sig_rx =-84;
13854: waveform_sig_rx =134;
13855: waveform_sig_rx =148;
13856: waveform_sig_rx =-153;
13857: waveform_sig_rx =160;
13858: waveform_sig_rx =144;
13859: waveform_sig_rx =-59;
13860: waveform_sig_rx =74;
13861: waveform_sig_rx =209;
13862: waveform_sig_rx =59;
13863: waveform_sig_rx =-23;
13864: waveform_sig_rx =243;
13865: waveform_sig_rx =151;
13866: waveform_sig_rx =-45;
13867: waveform_sig_rx =223;
13868: waveform_sig_rx =266;
13869: waveform_sig_rx =-64;
13870: waveform_sig_rx =263;
13871: waveform_sig_rx =82;
13872: waveform_sig_rx =185;
13873: waveform_sig_rx =171;
13874: waveform_sig_rx =240;
13875: waveform_sig_rx =81;
13876: waveform_sig_rx =259;
13877: waveform_sig_rx =310;
13878: waveform_sig_rx =10;
13879: waveform_sig_rx =404;
13880: waveform_sig_rx =232;
13881: waveform_sig_rx =73;
13882: waveform_sig_rx =370;
13883: waveform_sig_rx =321;
13884: waveform_sig_rx =59;
13885: waveform_sig_rx =362;
13886: waveform_sig_rx =365;
13887: waveform_sig_rx =90;
13888: waveform_sig_rx =322;
13889: waveform_sig_rx =378;
13890: waveform_sig_rx =186;
13891: waveform_sig_rx =191;
13892: waveform_sig_rx =510;
13893: waveform_sig_rx =229;
13894: waveform_sig_rx =203;
13895: waveform_sig_rx =444;
13896: waveform_sig_rx =374;
13897: waveform_sig_rx =191;
13898: waveform_sig_rx =453;
13899: waveform_sig_rx =406;
13900: waveform_sig_rx =288;
13901: waveform_sig_rx =313;
13902: waveform_sig_rx =526;
13903: waveform_sig_rx =341;
13904: waveform_sig_rx =222;
13905: waveform_sig_rx =605;
13906: waveform_sig_rx =391;
13907: waveform_sig_rx =242;
13908: waveform_sig_rx =563;
13909: waveform_sig_rx =490;
13910: waveform_sig_rx =265;
13911: waveform_sig_rx =551;
13912: waveform_sig_rx =345;
13913: waveform_sig_rx =519;
13914: waveform_sig_rx =418;
13915: waveform_sig_rx =490;
13916: waveform_sig_rx =371;
13917: waveform_sig_rx =511;
13918: waveform_sig_rx =564;
13919: waveform_sig_rx =310;
13920: waveform_sig_rx =630;
13921: waveform_sig_rx =522;
13922: waveform_sig_rx =319;
13923: waveform_sig_rx =639;
13924: waveform_sig_rx =609;
13925: waveform_sig_rx =302;
13926: waveform_sig_rx =674;
13927: waveform_sig_rx =664;
13928: waveform_sig_rx =350;
13929: waveform_sig_rx =632;
13930: waveform_sig_rx =680;
13931: waveform_sig_rx =421;
13932: waveform_sig_rx =505;
13933: waveform_sig_rx =759;
13934: waveform_sig_rx =469;
13935: waveform_sig_rx =514;
13936: waveform_sig_rx =686;
13937: waveform_sig_rx =642;
13938: waveform_sig_rx =477;
13939: waveform_sig_rx =669;
13940: waveform_sig_rx =710;
13941: waveform_sig_rx =516;
13942: waveform_sig_rx =583;
13943: waveform_sig_rx =843;
13944: waveform_sig_rx =543;
13945: waveform_sig_rx =522;
13946: waveform_sig_rx =874;
13947: waveform_sig_rx =588;
13948: waveform_sig_rx =538;
13949: waveform_sig_rx =800;
13950: waveform_sig_rx =714;
13951: waveform_sig_rx =563;
13952: waveform_sig_rx =797;
13953: waveform_sig_rx =595;
13954: waveform_sig_rx =798;
13955: waveform_sig_rx =634;
13956: waveform_sig_rx =756;
13957: waveform_sig_rx =615;
13958: waveform_sig_rx =712;
13959: waveform_sig_rx =834;
13960: waveform_sig_rx =533;
13961: waveform_sig_rx =852;
13962: waveform_sig_rx =807;
13963: waveform_sig_rx =544;
13964: waveform_sig_rx =930;
13965: waveform_sig_rx =844;
13966: waveform_sig_rx =501;
13967: waveform_sig_rx =978;
13968: waveform_sig_rx =845;
13969: waveform_sig_rx =582;
13970: waveform_sig_rx =919;
13971: waveform_sig_rx =862;
13972: waveform_sig_rx =674;
13973: waveform_sig_rx =764;
13974: waveform_sig_rx =967;
13975: waveform_sig_rx =742;
13976: waveform_sig_rx =767;
13977: waveform_sig_rx =908;
13978: waveform_sig_rx =910;
13979: waveform_sig_rx =686;
13980: waveform_sig_rx =908;
13981: waveform_sig_rx =969;
13982: waveform_sig_rx =681;
13983: waveform_sig_rx =813;
13984: waveform_sig_rx =1065;
13985: waveform_sig_rx =699;
13986: waveform_sig_rx =789;
13987: waveform_sig_rx =1057;
13988: waveform_sig_rx =769;
13989: waveform_sig_rx =809;
13990: waveform_sig_rx =982;
13991: waveform_sig_rx =939;
13992: waveform_sig_rx =803;
13993: waveform_sig_rx =951;
13994: waveform_sig_rx =841;
13995: waveform_sig_rx =980;
13996: waveform_sig_rx =817;
13997: waveform_sig_rx =1017;
13998: waveform_sig_rx =777;
13999: waveform_sig_rx =980;
14000: waveform_sig_rx =1050;
14001: waveform_sig_rx =701;
14002: waveform_sig_rx =1128;
14003: waveform_sig_rx =962;
14004: waveform_sig_rx =732;
14005: waveform_sig_rx =1184;
14006: waveform_sig_rx =987;
14007: waveform_sig_rx =722;
14008: waveform_sig_rx =1172;
14009: waveform_sig_rx =982;
14010: waveform_sig_rx =784;
14011: waveform_sig_rx =1122;
14012: waveform_sig_rx =1035;
14013: waveform_sig_rx =862;
14014: waveform_sig_rx =965;
14015: waveform_sig_rx =1116;
14016: waveform_sig_rx =925;
14017: waveform_sig_rx =889;
14018: waveform_sig_rx =1095;
14019: waveform_sig_rx =1089;
14020: waveform_sig_rx =781;
14021: waveform_sig_rx =1148;
14022: waveform_sig_rx =1097;
14023: waveform_sig_rx =831;
14024: waveform_sig_rx =1077;
14025: waveform_sig_rx =1171;
14026: waveform_sig_rx =889;
14027: waveform_sig_rx =989;
14028: waveform_sig_rx =1177;
14029: waveform_sig_rx =995;
14030: waveform_sig_rx =929;
14031: waveform_sig_rx =1138;
14032: waveform_sig_rx =1113;
14033: waveform_sig_rx =903;
14034: waveform_sig_rx =1144;
14035: waveform_sig_rx =1001;
14036: waveform_sig_rx =1113;
14037: waveform_sig_rx =1023;
14038: waveform_sig_rx =1188;
14039: waveform_sig_rx =895;
14040: waveform_sig_rx =1194;
14041: waveform_sig_rx =1132;
14042: waveform_sig_rx =848;
14043: waveform_sig_rx =1311;
14044: waveform_sig_rx =1039;
14045: waveform_sig_rx =909;
14046: waveform_sig_rx =1319;
14047: waveform_sig_rx =1050;
14048: waveform_sig_rx =892;
14049: waveform_sig_rx =1282;
14050: waveform_sig_rx =1076;
14051: waveform_sig_rx =967;
14052: waveform_sig_rx =1201;
14053: waveform_sig_rx =1167;
14054: waveform_sig_rx =994;
14055: waveform_sig_rx =1055;
14056: waveform_sig_rx =1272;
14057: waveform_sig_rx =1016;
14058: waveform_sig_rx =1006;
14059: waveform_sig_rx =1249;
14060: waveform_sig_rx =1159;
14061: waveform_sig_rx =920;
14062: waveform_sig_rx =1299;
14063: waveform_sig_rx =1153;
14064: waveform_sig_rx =984;
14065: waveform_sig_rx =1192;
14066: waveform_sig_rx =1217;
14067: waveform_sig_rx =1053;
14068: waveform_sig_rx =1041;
14069: waveform_sig_rx =1298;
14070: waveform_sig_rx =1108;
14071: waveform_sig_rx =992;
14072: waveform_sig_rx =1300;
14073: waveform_sig_rx =1165;
14074: waveform_sig_rx =976;
14075: waveform_sig_rx =1264;
14076: waveform_sig_rx =1029;
14077: waveform_sig_rx =1198;
14078: waveform_sig_rx =1085;
14079: waveform_sig_rx =1218;
14080: waveform_sig_rx =947;
14081: waveform_sig_rx =1274;
14082: waveform_sig_rx =1146;
14083: waveform_sig_rx =935;
14084: waveform_sig_rx =1403;
14085: waveform_sig_rx =1046;
14086: waveform_sig_rx =1028;
14087: waveform_sig_rx =1367;
14088: waveform_sig_rx =1088;
14089: waveform_sig_rx =1020;
14090: waveform_sig_rx =1292;
14091: waveform_sig_rx =1160;
14092: waveform_sig_rx =1028;
14093: waveform_sig_rx =1208;
14094: waveform_sig_rx =1280;
14095: waveform_sig_rx =951;
14096: waveform_sig_rx =1142;
14097: waveform_sig_rx =1333;
14098: waveform_sig_rx =1007;
14099: waveform_sig_rx =1116;
14100: waveform_sig_rx =1257;
14101: waveform_sig_rx =1154;
14102: waveform_sig_rx =997;
14103: waveform_sig_rx =1277;
14104: waveform_sig_rx =1183;
14105: waveform_sig_rx =1023;
14106: waveform_sig_rx =1201;
14107: waveform_sig_rx =1266;
14108: waveform_sig_rx =1070;
14109: waveform_sig_rx =1060;
14110: waveform_sig_rx =1322;
14111: waveform_sig_rx =1108;
14112: waveform_sig_rx =962;
14113: waveform_sig_rx =1353;
14114: waveform_sig_rx =1130;
14115: waveform_sig_rx =1001;
14116: waveform_sig_rx =1310;
14117: waveform_sig_rx =987;
14118: waveform_sig_rx =1267;
14119: waveform_sig_rx =1070;
14120: waveform_sig_rx =1197;
14121: waveform_sig_rx =998;
14122: waveform_sig_rx =1269;
14123: waveform_sig_rx =1124;
14124: waveform_sig_rx =970;
14125: waveform_sig_rx =1340;
14126: waveform_sig_rx =1066;
14127: waveform_sig_rx =1014;
14128: waveform_sig_rx =1319;
14129: waveform_sig_rx =1098;
14130: waveform_sig_rx =965;
14131: waveform_sig_rx =1280;
14132: waveform_sig_rx =1120;
14133: waveform_sig_rx =949;
14134: waveform_sig_rx =1206;
14135: waveform_sig_rx =1241;
14136: waveform_sig_rx =918;
14137: waveform_sig_rx =1160;
14138: waveform_sig_rx =1252;
14139: waveform_sig_rx =952;
14140: waveform_sig_rx =1098;
14141: waveform_sig_rx =1192;
14142: waveform_sig_rx =1124;
14143: waveform_sig_rx =972;
14144: waveform_sig_rx =1196;
14145: waveform_sig_rx =1156;
14146: waveform_sig_rx =949;
14147: waveform_sig_rx =1132;
14148: waveform_sig_rx =1239;
14149: waveform_sig_rx =948;
14150: waveform_sig_rx =1038;
14151: waveform_sig_rx =1311;
14152: waveform_sig_rx =1004;
14153: waveform_sig_rx =982;
14154: waveform_sig_rx =1305;
14155: waveform_sig_rx =1012;
14156: waveform_sig_rx =1020;
14157: waveform_sig_rx =1185;
14158: waveform_sig_rx =928;
14159: waveform_sig_rx =1240;
14160: waveform_sig_rx =954;
14161: waveform_sig_rx =1166;
14162: waveform_sig_rx =900;
14163: waveform_sig_rx =1170;
14164: waveform_sig_rx =1076;
14165: waveform_sig_rx =884;
14166: waveform_sig_rx =1260;
14167: waveform_sig_rx =988;
14168: waveform_sig_rx =896;
14169: waveform_sig_rx =1260;
14170: waveform_sig_rx =974;
14171: waveform_sig_rx =857;
14172: waveform_sig_rx =1223;
14173: waveform_sig_rx =1030;
14174: waveform_sig_rx =833;
14175: waveform_sig_rx =1157;
14176: waveform_sig_rx =1100;
14177: waveform_sig_rx =792;
14178: waveform_sig_rx =1113;
14179: waveform_sig_rx =1091;
14180: waveform_sig_rx =905;
14181: waveform_sig_rx =1003;
14182: waveform_sig_rx =1060;
14183: waveform_sig_rx =1062;
14184: waveform_sig_rx =822;
14185: waveform_sig_rx =1119;
14186: waveform_sig_rx =1066;
14187: waveform_sig_rx =784;
14188: waveform_sig_rx =1069;
14189: waveform_sig_rx =1124;
14190: waveform_sig_rx =781;
14191: waveform_sig_rx =983;
14192: waveform_sig_rx =1124;
14193: waveform_sig_rx =854;
14194: waveform_sig_rx =896;
14195: waveform_sig_rx =1098;
14196: waveform_sig_rx =923;
14197: waveform_sig_rx =876;
14198: waveform_sig_rx =1012;
14199: waveform_sig_rx =833;
14200: waveform_sig_rx =1043;
14201: waveform_sig_rx =838;
14202: waveform_sig_rx =1056;
14203: waveform_sig_rx =733;
14204: waveform_sig_rx =1072;
14205: waveform_sig_rx =910;
14206: waveform_sig_rx =731;
14207: waveform_sig_rx =1124;
14208: waveform_sig_rx =806;
14209: waveform_sig_rx =739;
14210: waveform_sig_rx =1103;
14211: waveform_sig_rx =814;
14212: waveform_sig_rx =663;
14213: waveform_sig_rx =1126;
14214: waveform_sig_rx =793;
14215: waveform_sig_rx =719;
14216: waveform_sig_rx =1046;
14217: waveform_sig_rx =853;
14218: waveform_sig_rx =726;
14219: waveform_sig_rx =919;
14220: waveform_sig_rx =926;
14221: waveform_sig_rx =799;
14222: waveform_sig_rx =748;
14223: waveform_sig_rx =955;
14224: waveform_sig_rx =852;
14225: waveform_sig_rx =599;
14226: waveform_sig_rx =1014;
14227: waveform_sig_rx =787;
14228: waveform_sig_rx =631;
14229: waveform_sig_rx =896;
14230: waveform_sig_rx =864;
14231: waveform_sig_rx =662;
14232: waveform_sig_rx =769;
14233: waveform_sig_rx =944;
14234: waveform_sig_rx =665;
14235: waveform_sig_rx =680;
14236: waveform_sig_rx =933;
14237: waveform_sig_rx =695;
14238: waveform_sig_rx =688;
14239: waveform_sig_rx =775;
14240: waveform_sig_rx =666;
14241: waveform_sig_rx =809;
14242: waveform_sig_rx =617;
14243: waveform_sig_rx =862;
14244: waveform_sig_rx =484;
14245: waveform_sig_rx =886;
14246: waveform_sig_rx =680;
14247: waveform_sig_rx =500;
14248: waveform_sig_rx =974;
14249: waveform_sig_rx =557;
14250: waveform_sig_rx =554;
14251: waveform_sig_rx =941;
14252: waveform_sig_rx =510;
14253: waveform_sig_rx =544;
14254: waveform_sig_rx =858;
14255: waveform_sig_rx =557;
14256: waveform_sig_rx =557;
14257: waveform_sig_rx =726;
14258: waveform_sig_rx =691;
14259: waveform_sig_rx =467;
14260: waveform_sig_rx =647;
14261: waveform_sig_rx =739;
14262: waveform_sig_rx =472;
14263: waveform_sig_rx =525;
14264: waveform_sig_rx =746;
14265: waveform_sig_rx =544;
14266: waveform_sig_rx =433;
14267: waveform_sig_rx =758;
14268: waveform_sig_rx =542;
14269: waveform_sig_rx =417;
14270: waveform_sig_rx =649;
14271: waveform_sig_rx =618;
14272: waveform_sig_rx =386;
14273: waveform_sig_rx =543;
14274: waveform_sig_rx =639;
14275: waveform_sig_rx =438;
14276: waveform_sig_rx =442;
14277: waveform_sig_rx =650;
14278: waveform_sig_rx =481;
14279: waveform_sig_rx =394;
14280: waveform_sig_rx =561;
14281: waveform_sig_rx =419;
14282: waveform_sig_rx =493;
14283: waveform_sig_rx =448;
14284: waveform_sig_rx =545;
14285: waveform_sig_rx =236;
14286: waveform_sig_rx =702;
14287: waveform_sig_rx =327;
14288: waveform_sig_rx =327;
14289: waveform_sig_rx =687;
14290: waveform_sig_rx =211;
14291: waveform_sig_rx =389;
14292: waveform_sig_rx =592;
14293: waveform_sig_rx =262;
14294: waveform_sig_rx =298;
14295: waveform_sig_rx =545;
14296: waveform_sig_rx =331;
14297: waveform_sig_rx =266;
14298: waveform_sig_rx =460;
14299: waveform_sig_rx =436;
14300: waveform_sig_rx =155;
14301: waveform_sig_rx =405;
14302: waveform_sig_rx =453;
14303: waveform_sig_rx =177;
14304: waveform_sig_rx =273;
14305: waveform_sig_rx =468;
14306: waveform_sig_rx =239;
14307: waveform_sig_rx =170;
14308: waveform_sig_rx =491;
14309: waveform_sig_rx =254;
14310: waveform_sig_rx =172;
14311: waveform_sig_rx =374;
14312: waveform_sig_rx =336;
14313: waveform_sig_rx =147;
14314: waveform_sig_rx =226;
14315: waveform_sig_rx =377;
14316: waveform_sig_rx =163;
14317: waveform_sig_rx =85;
14318: waveform_sig_rx =440;
14319: waveform_sig_rx =152;
14320: waveform_sig_rx =102;
14321: waveform_sig_rx =336;
14322: waveform_sig_rx =50;
14323: waveform_sig_rx =275;
14324: waveform_sig_rx =164;
14325: waveform_sig_rx =188;
14326: waveform_sig_rx =33;
14327: waveform_sig_rx =347;
14328: waveform_sig_rx =2;
14329: waveform_sig_rx =92;
14330: waveform_sig_rx =300;
14331: waveform_sig_rx =4;
14332: waveform_sig_rx =83;
14333: waveform_sig_rx =295;
14334: waveform_sig_rx =32;
14335: waveform_sig_rx =-19;
14336: waveform_sig_rx =300;
14337: waveform_sig_rx =0;
14338: waveform_sig_rx =-24;
14339: waveform_sig_rx =174;
14340: waveform_sig_rx =116;
14341: waveform_sig_rx =-158;
14342: waveform_sig_rx =129;
14343: waveform_sig_rx =163;
14344: waveform_sig_rx =-169;
14345: waveform_sig_rx =31;
14346: waveform_sig_rx =154;
14347: waveform_sig_rx =-96;
14348: waveform_sig_rx =-53;
14349: waveform_sig_rx =89;
14350: waveform_sig_rx =-32;
14351: waveform_sig_rx =-131;
14352: waveform_sig_rx =-3;
14353: waveform_sig_rx =129;
14354: waveform_sig_rx =-241;
14355: waveform_sig_rx =-34;
14356: waveform_sig_rx =131;
14357: waveform_sig_rx =-247;
14358: waveform_sig_rx =-111;
14359: waveform_sig_rx =127;
14360: waveform_sig_rx =-194;
14361: waveform_sig_rx =-106;
14362: waveform_sig_rx =-39;
14363: waveform_sig_rx =-204;
14364: waveform_sig_rx =-17;
14365: waveform_sig_rx =-189;
14366: waveform_sig_rx =-64;
14367: waveform_sig_rx =-256;
14368: waveform_sig_rx =33;
14369: waveform_sig_rx =-235;
14370: waveform_sig_rx =-219;
14371: waveform_sig_rx =2;
14372: waveform_sig_rx =-286;
14373: waveform_sig_rx =-272;
14374: waveform_sig_rx =4;
14375: waveform_sig_rx =-294;
14376: waveform_sig_rx =-375;
14377: waveform_sig_rx =44;
14378: waveform_sig_rx =-330;
14379: waveform_sig_rx =-358;
14380: waveform_sig_rx =-72;
14381: waveform_sig_rx =-230;
14382: waveform_sig_rx =-458;
14383: waveform_sig_rx =-136;
14384: waveform_sig_rx =-196;
14385: waveform_sig_rx =-418;
14386: waveform_sig_rx =-256;
14387: waveform_sig_rx =-189;
14388: waveform_sig_rx =-354;
14389: waveform_sig_rx =-379;
14390: waveform_sig_rx =-205;
14391: waveform_sig_rx =-286;
14392: waveform_sig_rx =-488;
14393: waveform_sig_rx =-260;
14394: waveform_sig_rx =-202;
14395: waveform_sig_rx =-587;
14396: waveform_sig_rx =-262;
14397: waveform_sig_rx =-218;
14398: waveform_sig_rx =-548;
14399: waveform_sig_rx =-359;
14400: waveform_sig_rx =-254;
14401: waveform_sig_rx =-485;
14402: waveform_sig_rx =-418;
14403: waveform_sig_rx =-406;
14404: waveform_sig_rx =-441;
14405: waveform_sig_rx =-342;
14406: waveform_sig_rx =-501;
14407: waveform_sig_rx =-343;
14408: waveform_sig_rx =-595;
14409: waveform_sig_rx =-270;
14410: waveform_sig_rx =-541;
14411: waveform_sig_rx =-565;
14412: waveform_sig_rx =-264;
14413: waveform_sig_rx =-591;
14414: waveform_sig_rx =-584;
14415: waveform_sig_rx =-243;
14416: waveform_sig_rx =-626;
14417: waveform_sig_rx =-643;
14418: waveform_sig_rx =-218;
14419: waveform_sig_rx =-676;
14420: waveform_sig_rx =-606;
14421: waveform_sig_rx =-344;
14422: waveform_sig_rx =-578;
14423: waveform_sig_rx =-701;
14424: waveform_sig_rx =-437;
14425: waveform_sig_rx =-505;
14426: waveform_sig_rx =-649;
14427: waveform_sig_rx =-586;
14428: waveform_sig_rx =-447;
14429: waveform_sig_rx =-620;
14430: waveform_sig_rx =-711;
14431: waveform_sig_rx =-424;
14432: waveform_sig_rx =-593;
14433: waveform_sig_rx =-793;
14434: waveform_sig_rx =-460;
14435: waveform_sig_rx =-531;
14436: waveform_sig_rx =-839;
14437: waveform_sig_rx =-516;
14438: waveform_sig_rx =-550;
14439: waveform_sig_rx =-773;
14440: waveform_sig_rx =-646;
14441: waveform_sig_rx =-538;
14442: waveform_sig_rx =-724;
14443: waveform_sig_rx =-685;
14444: waveform_sig_rx =-674;
14445: waveform_sig_rx =-686;
14446: waveform_sig_rx =-658;
14447: waveform_sig_rx =-732;
14448: waveform_sig_rx =-617;
14449: waveform_sig_rx =-887;
14450: waveform_sig_rx =-464;
14451: waveform_sig_rx =-852;
14452: waveform_sig_rx =-809;
14453: waveform_sig_rx =-499;
14454: waveform_sig_rx =-928;
14455: waveform_sig_rx =-794;
14456: waveform_sig_rx =-507;
14457: waveform_sig_rx =-958;
14458: waveform_sig_rx =-852;
14459: waveform_sig_rx =-518;
14460: waveform_sig_rx =-968;
14461: waveform_sig_rx =-800;
14462: waveform_sig_rx =-655;
14463: waveform_sig_rx =-821;
14464: waveform_sig_rx =-934;
14465: waveform_sig_rx =-698;
14466: waveform_sig_rx =-757;
14467: waveform_sig_rx =-916;
14468: waveform_sig_rx =-872;
14469: waveform_sig_rx =-635;
14470: waveform_sig_rx =-921;
14471: waveform_sig_rx =-957;
14472: waveform_sig_rx =-584;
14473: waveform_sig_rx =-929;
14474: waveform_sig_rx =-979;
14475: waveform_sig_rx =-664;
14476: waveform_sig_rx =-855;
14477: waveform_sig_rx =-990;
14478: waveform_sig_rx =-791;
14479: waveform_sig_rx =-793;
14480: waveform_sig_rx =-965;
14481: waveform_sig_rx =-934;
14482: waveform_sig_rx =-697;
14483: waveform_sig_rx =-981;
14484: waveform_sig_rx =-936;
14485: waveform_sig_rx =-842;
14486: waveform_sig_rx =-961;
14487: waveform_sig_rx =-879;
14488: waveform_sig_rx =-918;
14489: waveform_sig_rx =-886;
14490: waveform_sig_rx =-1099;
14491: waveform_sig_rx =-681;
14492: waveform_sig_rx =-1132;
14493: waveform_sig_rx =-988;
14494: waveform_sig_rx =-719;
14495: waveform_sig_rx =-1179;
14496: waveform_sig_rx =-944;
14497: waveform_sig_rx =-726;
14498: waveform_sig_rx =-1193;
14499: waveform_sig_rx =-945;
14500: waveform_sig_rx =-793;
14501: waveform_sig_rx =-1144;
14502: waveform_sig_rx =-973;
14503: waveform_sig_rx =-931;
14504: waveform_sig_rx =-952;
14505: waveform_sig_rx =-1171;
14506: waveform_sig_rx =-921;
14507: waveform_sig_rx =-902;
14508: waveform_sig_rx =-1163;
14509: waveform_sig_rx =-1009;
14510: waveform_sig_rx =-827;
14511: waveform_sig_rx =-1173;
14512: waveform_sig_rx =-1062;
14513: waveform_sig_rx =-858;
14514: waveform_sig_rx =-1110;
14515: waveform_sig_rx =-1105;
14516: waveform_sig_rx =-913;
14517: waveform_sig_rx =-991;
14518: waveform_sig_rx =-1182;
14519: waveform_sig_rx =-1001;
14520: waveform_sig_rx =-910;
14521: waveform_sig_rx =-1188;
14522: waveform_sig_rx =-1086;
14523: waveform_sig_rx =-857;
14524: waveform_sig_rx =-1198;
14525: waveform_sig_rx =-1048;
14526: waveform_sig_rx =-1016;
14527: waveform_sig_rx =-1112;
14528: waveform_sig_rx =-1038;
14529: waveform_sig_rx =-1064;
14530: waveform_sig_rx =-1075;
14531: waveform_sig_rx =-1208;
14532: waveform_sig_rx =-848;
14533: waveform_sig_rx =-1310;
14534: waveform_sig_rx =-1057;
14535: waveform_sig_rx =-928;
14536: waveform_sig_rx =-1321;
14537: waveform_sig_rx =-1016;
14538: waveform_sig_rx =-966;
14539: waveform_sig_rx =-1264;
14540: waveform_sig_rx =-1123;
14541: waveform_sig_rx =-950;
14542: waveform_sig_rx =-1199;
14543: waveform_sig_rx =-1198;
14544: waveform_sig_rx =-975;
14545: waveform_sig_rx =-1100;
14546: waveform_sig_rx =-1343;
14547: waveform_sig_rx =-926;
14548: waveform_sig_rx =-1104;
14549: waveform_sig_rx =-1278;
14550: waveform_sig_rx =-1087;
14551: waveform_sig_rx =-1001;
14552: waveform_sig_rx =-1233;
14553: waveform_sig_rx =-1173;
14554: waveform_sig_rx =-1001;
14555: waveform_sig_rx =-1202;
14556: waveform_sig_rx =-1240;
14557: waveform_sig_rx =-1014;
14558: waveform_sig_rx =-1093;
14559: waveform_sig_rx =-1303;
14560: waveform_sig_rx =-1084;
14561: waveform_sig_rx =-1017;
14562: waveform_sig_rx =-1323;
14563: waveform_sig_rx =-1165;
14564: waveform_sig_rx =-948;
14565: waveform_sig_rx =-1324;
14566: waveform_sig_rx =-1095;
14567: waveform_sig_rx =-1145;
14568: waveform_sig_rx =-1208;
14569: waveform_sig_rx =-1090;
14570: waveform_sig_rx =-1180;
14571: waveform_sig_rx =-1168;
14572: waveform_sig_rx =-1249;
14573: waveform_sig_rx =-958;
14574: waveform_sig_rx =-1344;
14575: waveform_sig_rx =-1095;
14576: waveform_sig_rx =-1033;
14577: waveform_sig_rx =-1309;
14578: waveform_sig_rx =-1136;
14579: waveform_sig_rx =-999;
14580: waveform_sig_rx =-1291;
14581: waveform_sig_rx =-1239;
14582: waveform_sig_rx =-935;
14583: waveform_sig_rx =-1310;
14584: waveform_sig_rx =-1234;
14585: waveform_sig_rx =-969;
14586: waveform_sig_rx =-1226;
14587: waveform_sig_rx =-1311;
14588: waveform_sig_rx =-945;
14589: waveform_sig_rx =-1187;
14590: waveform_sig_rx =-1226;
14591: waveform_sig_rx =-1152;
14592: waveform_sig_rx =-1038;
14593: waveform_sig_rx =-1270;
14594: waveform_sig_rx =-1202;
14595: waveform_sig_rx =-993;
14596: waveform_sig_rx =-1245;
14597: waveform_sig_rx =-1242;
14598: waveform_sig_rx =-1029;
14599: waveform_sig_rx =-1090;
14600: waveform_sig_rx =-1366;
14601: waveform_sig_rx =-1060;
14602: waveform_sig_rx =-1023;
14603: waveform_sig_rx =-1391;
14604: waveform_sig_rx =-1080;
14605: waveform_sig_rx =-1005;
14606: waveform_sig_rx =-1335;
14607: waveform_sig_rx =-1018;
14608: waveform_sig_rx =-1242;
14609: waveform_sig_rx =-1120;
14610: waveform_sig_rx =-1105;
14611: waveform_sig_rx =-1201;
14612: waveform_sig_rx =-1079;
14613: waveform_sig_rx =-1282;
14614: waveform_sig_rx =-953;
14615: waveform_sig_rx =-1305;
14616: waveform_sig_rx =-1150;
14617: waveform_sig_rx =-961;
14618: waveform_sig_rx =-1330;
14619: waveform_sig_rx =-1100;
14620: waveform_sig_rx =-935;
14621: waveform_sig_rx =-1313;
14622: waveform_sig_rx =-1131;
14623: waveform_sig_rx =-912;
14624: waveform_sig_rx =-1299;
14625: waveform_sig_rx =-1145;
14626: waveform_sig_rx =-942;
14627: waveform_sig_rx =-1212;
14628: waveform_sig_rx =-1238;
14629: waveform_sig_rx =-919;
14630: waveform_sig_rx =-1170;
14631: waveform_sig_rx =-1148;
14632: waveform_sig_rx =-1120;
14633: waveform_sig_rx =-973;
14634: waveform_sig_rx =-1200;
14635: waveform_sig_rx =-1180;
14636: waveform_sig_rx =-914;
14637: waveform_sig_rx =-1179;
14638: waveform_sig_rx =-1225;
14639: waveform_sig_rx =-897;
14640: waveform_sig_rx =-1085;
14641: waveform_sig_rx =-1262;
14642: waveform_sig_rx =-937;
14643: waveform_sig_rx =-1039;
14644: waveform_sig_rx =-1240;
14645: waveform_sig_rx =-1014;
14646: waveform_sig_rx =-967;
14647: waveform_sig_rx =-1192;
14648: waveform_sig_rx =-1017;
14649: waveform_sig_rx =-1143;
14650: waveform_sig_rx =-996;
14651: waveform_sig_rx =-1110;
14652: waveform_sig_rx =-1043;
14653: waveform_sig_rx =-1005;
14654: waveform_sig_rx =-1197;
14655: waveform_sig_rx =-783;
14656: waveform_sig_rx =-1255;
14657: waveform_sig_rx =-1017;
14658: waveform_sig_rx =-830;
14659: waveform_sig_rx =-1289;
14660: waveform_sig_rx =-937;
14661: waveform_sig_rx =-840;
14662: waveform_sig_rx =-1239;
14663: waveform_sig_rx =-994;
14664: waveform_sig_rx =-826;
14665: waveform_sig_rx =-1205;
14666: waveform_sig_rx =-977;
14667: waveform_sig_rx =-843;
14668: waveform_sig_rx =-1104;
14669: waveform_sig_rx =-1083;
14670: waveform_sig_rx =-844;
14671: waveform_sig_rx =-1012;
14672: waveform_sig_rx =-1024;
14673: waveform_sig_rx =-1018;
14674: waveform_sig_rx =-780;
14675: waveform_sig_rx =-1133;
14676: waveform_sig_rx =-1025;
14677: waveform_sig_rx =-726;
14678: waveform_sig_rx =-1132;
14679: waveform_sig_rx =-1011;
14680: waveform_sig_rx =-769;
14681: waveform_sig_rx =-1016;
14682: waveform_sig_rx =-1042;
14683: waveform_sig_rx =-846;
14684: waveform_sig_rx =-891;
14685: waveform_sig_rx =-1055;
14686: waveform_sig_rx =-899;
14687: waveform_sig_rx =-757;
14688: waveform_sig_rx =-1064;
14689: waveform_sig_rx =-849;
14690: waveform_sig_rx =-951;
14691: waveform_sig_rx =-865;
14692: waveform_sig_rx =-929;
14693: waveform_sig_rx =-830;
14694: waveform_sig_rx =-899;
14695: waveform_sig_rx =-977;
14696: waveform_sig_rx =-622;
14697: waveform_sig_rx =-1129;
14698: waveform_sig_rx =-790;
14699: waveform_sig_rx =-705;
14700: waveform_sig_rx =-1123;
14701: waveform_sig_rx =-724;
14702: waveform_sig_rx =-711;
14703: waveform_sig_rx =-1092;
14704: waveform_sig_rx =-732;
14705: waveform_sig_rx =-698;
14706: waveform_sig_rx =-1002;
14707: waveform_sig_rx =-777;
14708: waveform_sig_rx =-724;
14709: waveform_sig_rx =-850;
14710: waveform_sig_rx =-935;
14711: waveform_sig_rx =-656;
14712: waveform_sig_rx =-752;
14713: waveform_sig_rx =-916;
14714: waveform_sig_rx =-772;
14715: waveform_sig_rx =-617;
14716: waveform_sig_rx =-976;
14717: waveform_sig_rx =-727;
14718: waveform_sig_rx =-594;
14719: waveform_sig_rx =-902;
14720: waveform_sig_rx =-763;
14721: waveform_sig_rx =-607;
14722: waveform_sig_rx =-769;
14723: waveform_sig_rx =-859;
14724: waveform_sig_rx =-627;
14725: waveform_sig_rx =-657;
14726: waveform_sig_rx =-845;
14727: waveform_sig_rx =-686;
14728: waveform_sig_rx =-540;
14729: waveform_sig_rx =-860;
14730: waveform_sig_rx =-653;
14731: waveform_sig_rx =-692;
14732: waveform_sig_rx =-679;
14733: waveform_sig_rx =-681;
14734: waveform_sig_rx =-597;
14735: waveform_sig_rx =-760;
14736: waveform_sig_rx =-688;
14737: waveform_sig_rx =-459;
14738: waveform_sig_rx =-911;
14739: waveform_sig_rx =-482;
14740: waveform_sig_rx =-566;
14741: waveform_sig_rx =-836;
14742: waveform_sig_rx =-493;
14743: waveform_sig_rx =-534;
14744: waveform_sig_rx =-794;
14745: waveform_sig_rx =-553;
14746: waveform_sig_rx =-474;
14747: waveform_sig_rx =-752;
14748: waveform_sig_rx =-582;
14749: waveform_sig_rx =-457;
14750: waveform_sig_rx =-624;
14751: waveform_sig_rx =-713;
14752: waveform_sig_rx =-366;
14753: waveform_sig_rx =-584;
14754: waveform_sig_rx =-679;
14755: waveform_sig_rx =-462;
14756: waveform_sig_rx =-425;
14757: waveform_sig_rx =-699;
14758: waveform_sig_rx =-458;
14759: waveform_sig_rx =-409;
14760: waveform_sig_rx =-627;
14761: waveform_sig_rx =-536;
14762: waveform_sig_rx =-378;
14763: waveform_sig_rx =-483;
14764: waveform_sig_rx =-639;
14765: waveform_sig_rx =-348;
14766: waveform_sig_rx =-393;
14767: waveform_sig_rx =-629;
14768: waveform_sig_rx =-395;
14769: waveform_sig_rx =-288;
14770: waveform_sig_rx =-646;
14771: waveform_sig_rx =-322;
14772: waveform_sig_rx =-487;
14773: waveform_sig_rx =-458;
14774: waveform_sig_rx =-389;
14775: waveform_sig_rx =-393;
14776: waveform_sig_rx =-481;
14777: waveform_sig_rx =-382;
14778: waveform_sig_rx =-258;
14779: waveform_sig_rx =-585;
14780: waveform_sig_rx =-257;
14781: waveform_sig_rx =-317;
14782: waveform_sig_rx =-502;
14783: waveform_sig_rx =-271;
14784: waveform_sig_rx =-216;
14785: waveform_sig_rx =-538;
14786: waveform_sig_rx =-300;
14787: waveform_sig_rx =-152;
14788: waveform_sig_rx =-504;
14789: waveform_sig_rx =-283;
14790: waveform_sig_rx =-173;
14791: waveform_sig_rx =-387;
14792: waveform_sig_rx =-422;
14793: waveform_sig_rx =-75;
14794: waveform_sig_rx =-342;
14795: waveform_sig_rx =-385;
14796: waveform_sig_rx =-170;
14797: waveform_sig_rx =-171;
14798: waveform_sig_rx =-382;
14799: waveform_sig_rx =-176;
14800: waveform_sig_rx =-136;
14801: waveform_sig_rx =-292;
14802: waveform_sig_rx =-293;
14803: waveform_sig_rx =-47;
14804: waveform_sig_rx =-198;
14805: waveform_sig_rx =-387;
14806: waveform_sig_rx =6;
14807: waveform_sig_rx =-154;
14808: waveform_sig_rx =-363;
14809: waveform_sig_rx =-55;
14810: waveform_sig_rx =-61;
14811: waveform_sig_rx =-328;
14812: waveform_sig_rx =-28;
14813: waveform_sig_rx =-247;
14814: waveform_sig_rx =-78;
14815: waveform_sig_rx =-123;
14816: waveform_sig_rx =-107;
14817: waveform_sig_rx =-139;
14818: waveform_sig_rx =-128;
14819: waveform_sig_rx =36;
14820: waveform_sig_rx =-266;
14821: waveform_sig_rx =1;
14822: waveform_sig_rx =9;
14823: waveform_sig_rx =-259;
14824: waveform_sig_rx =20;
14825: waveform_sig_rx =82;
14826: waveform_sig_rx =-301;
14827: waveform_sig_rx =41;
14828: waveform_sig_rx =131;
14829: waveform_sig_rx =-245;
14830: waveform_sig_rx =38;
14831: waveform_sig_rx =119;
14832: waveform_sig_rx =-129;
14833: waveform_sig_rx =-78;
14834: waveform_sig_rx =218;
14835: waveform_sig_rx =-66;
14836: waveform_sig_rx =-29;
14837: waveform_sig_rx =98;
14838: waveform_sig_rx =137;
14839: waveform_sig_rx =-67;
14840: waveform_sig_rx =60;
14841: waveform_sig_rx =226;
14842: waveform_sig_rx =-29;
14843: waveform_sig_rx =-25;
14844: waveform_sig_rx =324;
14845: waveform_sig_rx =17;
14846: waveform_sig_rx =-44;
14847: waveform_sig_rx =307;
14848: waveform_sig_rx =67;
14849: waveform_sig_rx =5;
14850: waveform_sig_rx =216;
14851: waveform_sig_rx =215;
14852: waveform_sig_rx =0;
14853: waveform_sig_rx =225;
14854: waveform_sig_rx =53;
14855: waveform_sig_rx =232;
14856: waveform_sig_rx =112;
14857: waveform_sig_rx =219;
14858: waveform_sig_rx =129;
14859: waveform_sig_rx =137;
14860: waveform_sig_rx =361;
14861: waveform_sig_rx =-20;
14862: waveform_sig_rx =282;
14863: waveform_sig_rx =329;
14864: waveform_sig_rx =-14;
14865: waveform_sig_rx =377;
14866: waveform_sig_rx =378;
14867: waveform_sig_rx =-44;
14868: waveform_sig_rx =409;
14869: waveform_sig_rx =353;
14870: waveform_sig_rx =33;
14871: waveform_sig_rx =396;
14872: waveform_sig_rx =354;
14873: waveform_sig_rx =182;
14874: waveform_sig_rx =236;
14875: waveform_sig_rx =451;
14876: waveform_sig_rx =253;
14877: waveform_sig_rx =243;
14878: waveform_sig_rx =367;
14879: waveform_sig_rx =454;
14880: waveform_sig_rx =181;
14881: waveform_sig_rx =366;
14882: waveform_sig_rx =522;
14883: waveform_sig_rx =196;
14884: waveform_sig_rx =317;
14885: waveform_sig_rx =593;
14886: waveform_sig_rx =254;
14887: waveform_sig_rx =289;
14888: waveform_sig_rx =569;
14889: waveform_sig_rx =349;
14890: waveform_sig_rx =340;
14891: waveform_sig_rx =447;
14892: waveform_sig_rx =539;
14893: waveform_sig_rx =290;
14894: waveform_sig_rx =494;
14895: waveform_sig_rx =398;
14896: waveform_sig_rx =497;
14897: waveform_sig_rx =396;
14898: waveform_sig_rx =562;
14899: waveform_sig_rx =362;
14900: waveform_sig_rx =443;
14901: waveform_sig_rx =629;
14902: waveform_sig_rx =217;
14903: waveform_sig_rx =634;
14904: waveform_sig_rx =568;
14905: waveform_sig_rx =254;
14906: waveform_sig_rx =694;
14907: waveform_sig_rx =586;
14908: waveform_sig_rx =258;
14909: waveform_sig_rx =705;
14910: waveform_sig_rx =598;
14911: waveform_sig_rx =336;
14912: waveform_sig_rx =636;
14913: waveform_sig_rx =609;
14914: waveform_sig_rx =482;
14915: waveform_sig_rx =494;
14916: waveform_sig_rx =722;
14917: waveform_sig_rx =559;
14918: waveform_sig_rx =471;
14919: waveform_sig_rx =657;
14920: waveform_sig_rx =715;
14921: waveform_sig_rx =389;
14922: waveform_sig_rx =721;
14923: waveform_sig_rx =751;
14924: waveform_sig_rx =439;
14925: waveform_sig_rx =657;
14926: waveform_sig_rx =798;
14927: waveform_sig_rx =550;
14928: waveform_sig_rx =590;
14929: waveform_sig_rx =758;
14930: waveform_sig_rx =661;
14931: waveform_sig_rx =532;
14932: waveform_sig_rx =730;
14933: waveform_sig_rx =826;
14934: waveform_sig_rx =491;
14935: waveform_sig_rx =765;
14936: waveform_sig_rx =645;
14937: waveform_sig_rx =711;
14938: waveform_sig_rx =692;
14939: waveform_sig_rx =794;
14940: waveform_sig_rx =578;
14941: waveform_sig_rx =789;
14942: waveform_sig_rx =819;
14943: waveform_sig_rx =475;
14944: waveform_sig_rx =934;
14945: waveform_sig_rx =753;
14946: waveform_sig_rx =549;
14947: waveform_sig_rx =957;
14948: waveform_sig_rx =814;
14949: waveform_sig_rx =565;
14950: waveform_sig_rx =949;
14951: waveform_sig_rx =829;
14952: waveform_sig_rx =629;
14953: waveform_sig_rx =880;
14954: waveform_sig_rx =865;
14955: waveform_sig_rx =741;
14956: waveform_sig_rx =696;
14957: waveform_sig_rx =1011;
14958: waveform_sig_rx =768;
14959: waveform_sig_rx =658;
14960: waveform_sig_rx =990;
14961: waveform_sig_rx =902;
14962: waveform_sig_rx =618;
14963: waveform_sig_rx =988;
14964: waveform_sig_rx =869;
14965: waveform_sig_rx =733;
14966: waveform_sig_rx =855;
14967: waveform_sig_rx =958;
14968: waveform_sig_rx =832;
14969: waveform_sig_rx =731;
14970: waveform_sig_rx =1026;
14971: waveform_sig_rx =891;
14972: waveform_sig_rx =691;
14973: waveform_sig_rx =1022;
14974: waveform_sig_rx =965;
14975: waveform_sig_rx =704;
14976: waveform_sig_rx =1022;
14977: waveform_sig_rx =798;
14978: waveform_sig_rx =976;
14979: waveform_sig_rx =885;
14980: waveform_sig_rx =990;
14981: waveform_sig_rx =782;
14982: waveform_sig_rx =1001;
14983: waveform_sig_rx =1019;
14984: waveform_sig_rx =710;
14985: waveform_sig_rx =1132;
14986: waveform_sig_rx =901;
14987: waveform_sig_rx =773;
14988: waveform_sig_rx =1113;
14989: waveform_sig_rx =948;
14990: waveform_sig_rx =809;
14991: waveform_sig_rx =1063;
14992: waveform_sig_rx =1047;
14993: waveform_sig_rx =820;
14994: waveform_sig_rx =1003;
14995: waveform_sig_rx =1143;
14996: waveform_sig_rx =808;
14997: waveform_sig_rx =914;
14998: waveform_sig_rx =1206;
14999: waveform_sig_rx =827;
15000: waveform_sig_rx =948;
15001: waveform_sig_rx =1105;
15002: waveform_sig_rx =1028;
15003: waveform_sig_rx =866;
15004: waveform_sig_rx =1074;
15005: waveform_sig_rx =1098;
15006: waveform_sig_rx =884;
15007: waveform_sig_rx =999;
15008: waveform_sig_rx =1172;
15009: waveform_sig_rx =938;
15010: waveform_sig_rx =917;
15011: waveform_sig_rx =1211;
15012: waveform_sig_rx =1014;
15013: waveform_sig_rx =874;
15014: waveform_sig_rx =1209;
15015: waveform_sig_rx =1077;
15016: waveform_sig_rx =883;
15017: waveform_sig_rx =1204;
15018: waveform_sig_rx =914;
15019: waveform_sig_rx =1140;
15020: waveform_sig_rx =1023;
15021: waveform_sig_rx =1124;
15022: waveform_sig_rx =957;
15023: waveform_sig_rx =1147;
15024: waveform_sig_rx =1116;
15025: waveform_sig_rx =900;
15026: waveform_sig_rx =1250;
15027: waveform_sig_rx =1046;
15028: waveform_sig_rx =961;
15029: waveform_sig_rx =1224;
15030: waveform_sig_rx =1150;
15031: waveform_sig_rx =865;
15032: waveform_sig_rx =1209;
15033: waveform_sig_rx =1194;
15034: waveform_sig_rx =849;
15035: waveform_sig_rx =1218;
15036: waveform_sig_rx =1223;
15037: waveform_sig_rx =870;
15038: waveform_sig_rx =1138;
15039: waveform_sig_rx =1235;
15040: waveform_sig_rx =1004;
15041: waveform_sig_rx =1069;
15042: waveform_sig_rx =1140;
15043: waveform_sig_rx =1209;
15044: waveform_sig_rx =924;
15045: waveform_sig_rx =1221;
15046: waveform_sig_rx =1205;
15047: waveform_sig_rx =952;
15048: waveform_sig_rx =1137;
15049: waveform_sig_rx =1271;
15050: waveform_sig_rx =1034;
15051: waveform_sig_rx =1012;
15052: waveform_sig_rx =1326;
15053: waveform_sig_rx =1059;
15054: waveform_sig_rx =964;
15055: waveform_sig_rx =1350;
15056: waveform_sig_rx =1095;
15057: waveform_sig_rx =1037;
15058: waveform_sig_rx =1269;
15059: waveform_sig_rx =975;
15060: waveform_sig_rx =1311;
15061: waveform_sig_rx =1013;
15062: waveform_sig_rx =1223;
15063: waveform_sig_rx =1047;
15064: waveform_sig_rx =1148;
15065: waveform_sig_rx =1243;
15066: waveform_sig_rx =934;
15067: waveform_sig_rx =1275;
15068: waveform_sig_rx =1166;
15069: waveform_sig_rx =909;
15070: waveform_sig_rx =1362;
15071: waveform_sig_rx =1151;
15072: waveform_sig_rx =897;
15073: waveform_sig_rx =1358;
15074: waveform_sig_rx =1145;
15075: waveform_sig_rx =942;
15076: waveform_sig_rx =1291;
15077: waveform_sig_rx =1207;
15078: waveform_sig_rx =982;
15079: waveform_sig_rx =1184;
15080: waveform_sig_rx =1270;
15081: waveform_sig_rx =1073;
15082: waveform_sig_rx =1092;
15083: waveform_sig_rx =1227;
15084: waveform_sig_rx =1235;
15085: waveform_sig_rx =949;
15086: waveform_sig_rx =1270;
15087: waveform_sig_rx =1253;
15088: waveform_sig_rx =978;
15089: waveform_sig_rx =1205;
15090: waveform_sig_rx =1320;
15091: waveform_sig_rx =996;
15092: waveform_sig_rx =1076;
15093: waveform_sig_rx =1340;
15094: waveform_sig_rx =1037;
15095: waveform_sig_rx =1075;
15096: waveform_sig_rx =1282;
15097: waveform_sig_rx =1134;
15098: waveform_sig_rx =1090;
15099: waveform_sig_rx =1183;
15100: waveform_sig_rx =1072;
15101: waveform_sig_rx =1263;
15102: waveform_sig_rx =1025;
15103: waveform_sig_rx =1302;
15104: waveform_sig_rx =951;
15105: waveform_sig_rx =1236;
15106: waveform_sig_rx =1211;
15107: waveform_sig_rx =878;
15108: waveform_sig_rx =1368;
15109: waveform_sig_rx =1070;
15110: waveform_sig_rx =934;
15111: waveform_sig_rx =1354;
15112: waveform_sig_rx =1085;
15113: waveform_sig_rx =933;
15114: waveform_sig_rx =1317;
15115: waveform_sig_rx =1127;
15116: waveform_sig_rx =956;
15117: waveform_sig_rx =1257;
15118: waveform_sig_rx =1167;
15119: waveform_sig_rx =967;
15120: waveform_sig_rx =1137;
15121: waveform_sig_rx =1209;
15122: waveform_sig_rx =1069;
15123: waveform_sig_rx =1019;
15124: waveform_sig_rx =1207;
15125: waveform_sig_rx =1196;
15126: waveform_sig_rx =868;
15127: waveform_sig_rx =1299;
15128: waveform_sig_rx =1130;
15129: waveform_sig_rx =910;
15130: waveform_sig_rx =1217;
15131: waveform_sig_rx =1172;
15132: waveform_sig_rx =974;
15133: waveform_sig_rx =1069;
15134: waveform_sig_rx =1218;
15135: waveform_sig_rx =1047;
15136: waveform_sig_rx =981;
15137: waveform_sig_rx =1205;
15138: waveform_sig_rx =1122;
15139: waveform_sig_rx =942;
15140: waveform_sig_rx =1161;
15141: waveform_sig_rx =1003;
15142: waveform_sig_rx =1117;
15143: waveform_sig_rx =1011;
15144: waveform_sig_rx =1189;
15145: waveform_sig_rx =851;
15146: waveform_sig_rx =1232;
15147: waveform_sig_rx =1058;
15148: waveform_sig_rx =848;
15149: waveform_sig_rx =1324;
15150: waveform_sig_rx =934;
15151: waveform_sig_rx =931;
15152: waveform_sig_rx =1282;
15153: waveform_sig_rx =951;
15154: waveform_sig_rx =883;
15155: waveform_sig_rx =1214;
15156: waveform_sig_rx =980;
15157: waveform_sig_rx =904;
15158: waveform_sig_rx =1126;
15159: waveform_sig_rx =1088;
15160: waveform_sig_rx =899;
15161: waveform_sig_rx =995;
15162: waveform_sig_rx =1155;
15163: waveform_sig_rx =925;
15164: waveform_sig_rx =890;
15165: waveform_sig_rx =1186;
15166: waveform_sig_rx =989;
15167: waveform_sig_rx =801;
15168: waveform_sig_rx =1211;
15169: waveform_sig_rx =961;
15170: waveform_sig_rx =870;
15171: waveform_sig_rx =1055;
15172: waveform_sig_rx =1059;
15173: waveform_sig_rx =909;
15174: waveform_sig_rx =892;
15175: waveform_sig_rx =1136;
15176: waveform_sig_rx =911;
15177: waveform_sig_rx =794;
15178: waveform_sig_rx =1142;
15179: waveform_sig_rx =944;
15180: waveform_sig_rx =803;
15181: waveform_sig_rx =1076;
15182: waveform_sig_rx =836;
15183: waveform_sig_rx =1004;
15184: waveform_sig_rx =906;
15185: waveform_sig_rx =988;
15186: waveform_sig_rx =745;
15187: waveform_sig_rx =1106;
15188: waveform_sig_rx =839;
15189: waveform_sig_rx =785;
15190: waveform_sig_rx =1132;
15191: waveform_sig_rx =757;
15192: waveform_sig_rx =819;
15193: waveform_sig_rx =1055;
15194: waveform_sig_rx =801;
15195: waveform_sig_rx =745;
15196: waveform_sig_rx =1013;
15197: waveform_sig_rx =870;
15198: waveform_sig_rx =707;
15199: waveform_sig_rx =929;
15200: waveform_sig_rx =959;
15201: waveform_sig_rx =650;
15202: waveform_sig_rx =863;
15203: waveform_sig_rx =992;
15204: waveform_sig_rx =670;
15205: waveform_sig_rx =775;
15206: waveform_sig_rx =951;
15207: waveform_sig_rx =764;
15208: waveform_sig_rx =676;
15209: waveform_sig_rx =947;
15210: waveform_sig_rx =780;
15211: waveform_sig_rx =696;
15212: waveform_sig_rx =825;
15213: waveform_sig_rx =895;
15214: waveform_sig_rx =672;
15215: waveform_sig_rx =691;
15216: waveform_sig_rx =971;
15217: waveform_sig_rx =672;
15218: waveform_sig_rx =617;
15219: waveform_sig_rx =979;
15220: waveform_sig_rx =670;
15221: waveform_sig_rx =650;
15222: waveform_sig_rx =890;
15223: waveform_sig_rx =574;
15224: waveform_sig_rx =865;
15225: waveform_sig_rx =660;
15226: waveform_sig_rx =766;
15227: waveform_sig_rx =571;
15228: waveform_sig_rx =831;
15229: waveform_sig_rx =650;
15230: waveform_sig_rx =591;
15231: waveform_sig_rx =853;
15232: waveform_sig_rx =601;
15233: waveform_sig_rx =574;
15234: waveform_sig_rx =848;
15235: waveform_sig_rx =646;
15236: waveform_sig_rx =474;
15237: waveform_sig_rx =857;
15238: waveform_sig_rx =630;
15239: waveform_sig_rx =492;
15240: waveform_sig_rx =776;
15241: waveform_sig_rx =711;
15242: waveform_sig_rx =406;
15243: waveform_sig_rx =705;
15244: waveform_sig_rx =743;
15245: waveform_sig_rx =446;
15246: waveform_sig_rx =607;
15247: waveform_sig_rx =688;
15248: waveform_sig_rx =559;
15249: waveform_sig_rx =491;
15250: waveform_sig_rx =661;
15251: waveform_sig_rx =630;
15252: waveform_sig_rx =427;
15253: waveform_sig_rx =567;
15254: waveform_sig_rx =740;
15255: waveform_sig_rx =345;
15256: waveform_sig_rx =517;
15257: waveform_sig_rx =727;
15258: waveform_sig_rx =353;
15259: waveform_sig_rx =473;
15260: waveform_sig_rx =690;
15261: waveform_sig_rx =405;
15262: waveform_sig_rx =459;
15263: waveform_sig_rx =545;
15264: waveform_sig_rx =358;
15265: waveform_sig_rx =619;
15266: waveform_sig_rx =372;
15267: waveform_sig_rx =545;
15268: waveform_sig_rx =313;
15269: waveform_sig_rx =561;
15270: waveform_sig_rx =430;
15271: waveform_sig_rx =292;
15272: waveform_sig_rx =594;
15273: waveform_sig_rx =389;
15274: waveform_sig_rx =255;
15275: waveform_sig_rx =622;
15276: waveform_sig_rx =347;
15277: waveform_sig_rx =163;
15278: waveform_sig_rx =658;
15279: waveform_sig_rx =287;
15280: waveform_sig_rx =226;
15281: waveform_sig_rx =537;
15282: waveform_sig_rx =371;
15283: waveform_sig_rx =160;
15284: waveform_sig_rx =428;
15285: waveform_sig_rx =400;
15286: waveform_sig_rx =209;
15287: waveform_sig_rx =310;
15288: waveform_sig_rx =373;
15289: waveform_sig_rx =322;
15290: waveform_sig_rx =148;
15291: waveform_sig_rx =412;
15292: waveform_sig_rx =354;
15293: waveform_sig_rx =95;
15294: waveform_sig_rx =375;
15295: waveform_sig_rx =415;
15296: waveform_sig_rx =28;
15297: waveform_sig_rx =343;
15298: waveform_sig_rx =378;
15299: waveform_sig_rx =87;
15300: waveform_sig_rx =239;
15301: waveform_sig_rx =343;
15302: waveform_sig_rx =184;
15303: waveform_sig_rx =145;
15304: waveform_sig_rx =244;
15305: waveform_sig_rx =119;
15306: waveform_sig_rx =261;
15307: waveform_sig_rx =90;
15308: waveform_sig_rx =267;
15309: waveform_sig_rx =-2;
15310: waveform_sig_rx =306;
15311: waveform_sig_rx =120;
15312: waveform_sig_rx =-19;
15313: waveform_sig_rx =343;
15314: waveform_sig_rx =52;
15315: waveform_sig_rx =-42;
15316: waveform_sig_rx =412;
15317: waveform_sig_rx =-6;
15318: waveform_sig_rx =-88;
15319: waveform_sig_rx =392;
15320: waveform_sig_rx =-97;
15321: waveform_sig_rx =-12;
15322: waveform_sig_rx =222;
15323: waveform_sig_rx =30;
15324: waveform_sig_rx =-54;
15325: waveform_sig_rx =89;
15326: waveform_sig_rx =116;
15327: waveform_sig_rx =-53;
15328: waveform_sig_rx =-52;
15329: waveform_sig_rx =152;
15330: waveform_sig_rx =-22;
15331: waveform_sig_rx =-164;
15332: waveform_sig_rx =172;
15333: waveform_sig_rx =-16;
15334: waveform_sig_rx =-210;
15335: waveform_sig_rx =87;
15336: waveform_sig_rx =38;
15337: waveform_sig_rx =-228;
15338: waveform_sig_rx =9;
15339: waveform_sig_rx =15;
15340: waveform_sig_rx =-173;
15341: waveform_sig_rx =-131;
15342: waveform_sig_rx =39;
15343: waveform_sig_rx =-98;
15344: waveform_sig_rx =-192;
15345: waveform_sig_rx =-56;
15346: waveform_sig_rx =-132;
15347: waveform_sig_rx =-68;
15348: waveform_sig_rx =-177;
15349: waveform_sig_rx =-33;
15350: waveform_sig_rx =-357;
15351: waveform_sig_rx =62;
15352: waveform_sig_rx =-263;
15353: waveform_sig_rx =-332;
15354: waveform_sig_rx =79;
15355: waveform_sig_rx =-371;
15356: waveform_sig_rx =-287;
15357: waveform_sig_rx =48;
15358: waveform_sig_rx =-398;
15359: waveform_sig_rx =-298;
15360: waveform_sig_rx =19;
15361: waveform_sig_rx =-371;
15362: waveform_sig_rx =-266;
15363: waveform_sig_rx =-148;
15364: waveform_sig_rx =-217;
15365: waveform_sig_rx =-399;
15366: waveform_sig_rx =-231;
15367: waveform_sig_rx =-144;
15368: waveform_sig_rx =-404;
15369: waveform_sig_rx =-346;
15370: waveform_sig_rx =-105;
15371: waveform_sig_rx =-385;
15372: waveform_sig_rx =-441;
15373: waveform_sig_rx =-96;
15374: waveform_sig_rx =-375;
15375: waveform_sig_rx =-473;
15376: waveform_sig_rx =-204;
15377: waveform_sig_rx =-290;
15378: waveform_sig_rx =-476;
15379: waveform_sig_rx =-333;
15380: waveform_sig_rx =-259;
15381: waveform_sig_rx =-447;
15382: waveform_sig_rx =-473;
15383: waveform_sig_rx =-190;
15384: waveform_sig_rx =-457;
15385: waveform_sig_rx =-492;
15386: waveform_sig_rx =-311;
15387: waveform_sig_rx =-496;
15388: waveform_sig_rx =-357;
15389: waveform_sig_rx =-437;
15390: waveform_sig_rx =-396;
15391: waveform_sig_rx =-609;
15392: waveform_sig_rx =-225;
15393: waveform_sig_rx =-599;
15394: waveform_sig_rx =-543;
15395: waveform_sig_rx =-243;
15396: waveform_sig_rx =-656;
15397: waveform_sig_rx =-517;
15398: waveform_sig_rx =-293;
15399: waveform_sig_rx =-671;
15400: waveform_sig_rx =-570;
15401: waveform_sig_rx =-320;
15402: waveform_sig_rx =-628;
15403: waveform_sig_rx =-584;
15404: waveform_sig_rx =-461;
15405: waveform_sig_rx =-476;
15406: waveform_sig_rx =-740;
15407: waveform_sig_rx =-471;
15408: waveform_sig_rx =-439;
15409: waveform_sig_rx =-750;
15410: waveform_sig_rx =-586;
15411: waveform_sig_rx =-411;
15412: waveform_sig_rx =-698;
15413: waveform_sig_rx =-678;
15414: waveform_sig_rx =-435;
15415: waveform_sig_rx =-667;
15416: waveform_sig_rx =-716;
15417: waveform_sig_rx =-563;
15418: waveform_sig_rx =-538;
15419: waveform_sig_rx =-767;
15420: waveform_sig_rx =-648;
15421: waveform_sig_rx =-453;
15422: waveform_sig_rx =-802;
15423: waveform_sig_rx =-733;
15424: waveform_sig_rx =-430;
15425: waveform_sig_rx =-808;
15426: waveform_sig_rx =-703;
15427: waveform_sig_rx =-614;
15428: waveform_sig_rx =-794;
15429: waveform_sig_rx =-580;
15430: waveform_sig_rx =-748;
15431: waveform_sig_rx =-661;
15432: waveform_sig_rx =-845;
15433: waveform_sig_rx =-518;
15434: waveform_sig_rx =-868;
15435: waveform_sig_rx =-791;
15436: waveform_sig_rx =-548;
15437: waveform_sig_rx =-925;
15438: waveform_sig_rx =-775;
15439: waveform_sig_rx =-584;
15440: waveform_sig_rx =-883;
15441: waveform_sig_rx =-870;
15442: waveform_sig_rx =-585;
15443: waveform_sig_rx =-862;
15444: waveform_sig_rx =-899;
15445: waveform_sig_rx =-641;
15446: waveform_sig_rx =-738;
15447: waveform_sig_rx =-1050;
15448: waveform_sig_rx =-628;
15449: waveform_sig_rx =-766;
15450: waveform_sig_rx =-988;
15451: waveform_sig_rx =-766;
15452: waveform_sig_rx =-735;
15453: waveform_sig_rx =-897;
15454: waveform_sig_rx =-909;
15455: waveform_sig_rx =-728;
15456: waveform_sig_rx =-840;
15457: waveform_sig_rx =-1009;
15458: waveform_sig_rx =-756;
15459: waveform_sig_rx =-760;
15460: waveform_sig_rx =-1063;
15461: waveform_sig_rx =-827;
15462: waveform_sig_rx =-735;
15463: waveform_sig_rx =-1051;
15464: waveform_sig_rx =-920;
15465: waveform_sig_rx =-701;
15466: waveform_sig_rx =-1034;
15467: waveform_sig_rx =-884;
15468: waveform_sig_rx =-852;
15469: waveform_sig_rx =-990;
15470: waveform_sig_rx =-826;
15471: waveform_sig_rx =-977;
15472: waveform_sig_rx =-868;
15473: waveform_sig_rx =-1062;
15474: waveform_sig_rx =-760;
15475: waveform_sig_rx =-1063;
15476: waveform_sig_rx =-970;
15477: waveform_sig_rx =-800;
15478: waveform_sig_rx =-1062;
15479: waveform_sig_rx =-1014;
15480: waveform_sig_rx =-770;
15481: waveform_sig_rx =-1070;
15482: waveform_sig_rx =-1125;
15483: waveform_sig_rx =-703;
15484: waveform_sig_rx =-1123;
15485: waveform_sig_rx =-1097;
15486: waveform_sig_rx =-781;
15487: waveform_sig_rx =-1049;
15488: waveform_sig_rx =-1159;
15489: waveform_sig_rx =-849;
15490: waveform_sig_rx =-1017;
15491: waveform_sig_rx =-1077;
15492: waveform_sig_rx =-1064;
15493: waveform_sig_rx =-880;
15494: waveform_sig_rx =-1092;
15495: waveform_sig_rx =-1157;
15496: waveform_sig_rx =-845;
15497: waveform_sig_rx =-1082;
15498: waveform_sig_rx =-1181;
15499: waveform_sig_rx =-927;
15500: waveform_sig_rx =-977;
15501: waveform_sig_rx =-1252;
15502: waveform_sig_rx =-996;
15503: waveform_sig_rx =-903;
15504: waveform_sig_rx =-1257;
15505: waveform_sig_rx =-1029;
15506: waveform_sig_rx =-911;
15507: waveform_sig_rx =-1212;
15508: waveform_sig_rx =-986;
15509: waveform_sig_rx =-1124;
15510: waveform_sig_rx =-1084;
15511: waveform_sig_rx =-1015;
15512: waveform_sig_rx =-1169;
15513: waveform_sig_rx =-972;
15514: waveform_sig_rx =-1279;
15515: waveform_sig_rx =-897;
15516: waveform_sig_rx =-1190;
15517: waveform_sig_rx =-1191;
15518: waveform_sig_rx =-861;
15519: waveform_sig_rx =-1270;
15520: waveform_sig_rx =-1171;
15521: waveform_sig_rx =-829;
15522: waveform_sig_rx =-1319;
15523: waveform_sig_rx =-1174;
15524: waveform_sig_rx =-861;
15525: waveform_sig_rx =-1326;
15526: waveform_sig_rx =-1136;
15527: waveform_sig_rx =-962;
15528: waveform_sig_rx =-1169;
15529: waveform_sig_rx =-1256;
15530: waveform_sig_rx =-1009;
15531: waveform_sig_rx =-1101;
15532: waveform_sig_rx =-1216;
15533: waveform_sig_rx =-1177;
15534: waveform_sig_rx =-958;
15535: waveform_sig_rx =-1241;
15536: waveform_sig_rx =-1221;
15537: waveform_sig_rx =-943;
15538: waveform_sig_rx =-1217;
15539: waveform_sig_rx =-1250;
15540: waveform_sig_rx =-983;
15541: waveform_sig_rx =-1091;
15542: waveform_sig_rx =-1339;
15543: waveform_sig_rx =-1030;
15544: waveform_sig_rx =-1066;
15545: waveform_sig_rx =-1323;
15546: waveform_sig_rx =-1102;
15547: waveform_sig_rx =-1043;
15548: waveform_sig_rx =-1234;
15549: waveform_sig_rx =-1140;
15550: waveform_sig_rx =-1199;
15551: waveform_sig_rx =-1093;
15552: waveform_sig_rx =-1184;
15553: waveform_sig_rx =-1159;
15554: waveform_sig_rx =-1082;
15555: waveform_sig_rx =-1381;
15556: waveform_sig_rx =-882;
15557: waveform_sig_rx =-1375;
15558: waveform_sig_rx =-1185;
15559: waveform_sig_rx =-912;
15560: waveform_sig_rx =-1424;
15561: waveform_sig_rx =-1104;
15562: waveform_sig_rx =-979;
15563: waveform_sig_rx =-1350;
15564: waveform_sig_rx =-1174;
15565: waveform_sig_rx =-985;
15566: waveform_sig_rx =-1308;
15567: waveform_sig_rx =-1204;
15568: waveform_sig_rx =-1009;
15569: waveform_sig_rx =-1195;
15570: waveform_sig_rx =-1297;
15571: waveform_sig_rx =-1024;
15572: waveform_sig_rx =-1157;
15573: waveform_sig_rx =-1232;
15574: waveform_sig_rx =-1217;
15575: waveform_sig_rx =-955;
15576: waveform_sig_rx =-1263;
15577: waveform_sig_rx =-1242;
15578: waveform_sig_rx =-905;
15579: waveform_sig_rx =-1305;
15580: waveform_sig_rx =-1233;
15581: waveform_sig_rx =-988;
15582: waveform_sig_rx =-1194;
15583: waveform_sig_rx =-1245;
15584: waveform_sig_rx =-1114;
15585: waveform_sig_rx =-1073;
15586: waveform_sig_rx =-1250;
15587: waveform_sig_rx =-1215;
15588: waveform_sig_rx =-942;
15589: waveform_sig_rx =-1294;
15590: waveform_sig_rx =-1168;
15591: waveform_sig_rx =-1128;
15592: waveform_sig_rx =-1173;
15593: waveform_sig_rx =-1111;
15594: waveform_sig_rx =-1124;
15595: waveform_sig_rx =-1153;
15596: waveform_sig_rx =-1261;
15597: waveform_sig_rx =-898;
15598: waveform_sig_rx =-1352;
15599: waveform_sig_rx =-1072;
15600: waveform_sig_rx =-975;
15601: waveform_sig_rx =-1361;
15602: waveform_sig_rx =-1055;
15603: waveform_sig_rx =-966;
15604: waveform_sig_rx =-1313;
15605: waveform_sig_rx =-1107;
15606: waveform_sig_rx =-942;
15607: waveform_sig_rx =-1272;
15608: waveform_sig_rx =-1108;
15609: waveform_sig_rx =-1006;
15610: waveform_sig_rx =-1121;
15611: waveform_sig_rx =-1271;
15612: waveform_sig_rx =-998;
15613: waveform_sig_rx =-1068;
15614: waveform_sig_rx =-1254;
15615: waveform_sig_rx =-1117;
15616: waveform_sig_rx =-913;
15617: waveform_sig_rx =-1307;
15618: waveform_sig_rx =-1092;
15619: waveform_sig_rx =-925;
15620: waveform_sig_rx =-1225;
15621: waveform_sig_rx =-1121;
15622: waveform_sig_rx =-1014;
15623: waveform_sig_rx =-1051;
15624: waveform_sig_rx =-1241;
15625: waveform_sig_rx =-1045;
15626: waveform_sig_rx =-932;
15627: waveform_sig_rx =-1268;
15628: waveform_sig_rx =-1068;
15629: waveform_sig_rx =-860;
15630: waveform_sig_rx =-1263;
15631: waveform_sig_rx =-994;
15632: waveform_sig_rx =-1084;
15633: waveform_sig_rx =-1096;
15634: waveform_sig_rx =-1012;
15635: waveform_sig_rx =-1061;
15636: waveform_sig_rx =-1065;
15637: waveform_sig_rx =-1128;
15638: waveform_sig_rx =-843;
15639: waveform_sig_rx =-1258;
15640: waveform_sig_rx =-982;
15641: waveform_sig_rx =-915;
15642: waveform_sig_rx =-1230;
15643: waveform_sig_rx =-952;
15644: waveform_sig_rx =-892;
15645: waveform_sig_rx =-1180;
15646: waveform_sig_rx =-1011;
15647: waveform_sig_rx =-850;
15648: waveform_sig_rx =-1146;
15649: waveform_sig_rx =-1037;
15650: waveform_sig_rx =-874;
15651: waveform_sig_rx =-992;
15652: waveform_sig_rx =-1192;
15653: waveform_sig_rx =-796;
15654: waveform_sig_rx =-969;
15655: waveform_sig_rx =-1132;
15656: waveform_sig_rx =-906;
15657: waveform_sig_rx =-880;
15658: waveform_sig_rx =-1106;
15659: waveform_sig_rx =-938;
15660: waveform_sig_rx =-863;
15661: waveform_sig_rx =-1000;
15662: waveform_sig_rx =-1057;
15663: waveform_sig_rx =-836;
15664: waveform_sig_rx =-882;
15665: waveform_sig_rx =-1158;
15666: waveform_sig_rx =-815;
15667: waveform_sig_rx =-839;
15668: waveform_sig_rx =-1127;
15669: waveform_sig_rx =-861;
15670: waveform_sig_rx =-774;
15671: waveform_sig_rx =-1086;
15672: waveform_sig_rx =-814;
15673: waveform_sig_rx =-944;
15674: waveform_sig_rx =-905;
15675: waveform_sig_rx =-831;
15676: waveform_sig_rx =-909;
15677: waveform_sig_rx =-873;
15678: waveform_sig_rx =-934;
15679: waveform_sig_rx =-698;
15680: waveform_sig_rx =-1042;
15681: waveform_sig_rx =-808;
15682: waveform_sig_rx =-733;
15683: waveform_sig_rx =-1008;
15684: waveform_sig_rx =-825;
15685: waveform_sig_rx =-676;
15686: waveform_sig_rx =-1027;
15687: waveform_sig_rx =-856;
15688: waveform_sig_rx =-603;
15689: waveform_sig_rx =-1021;
15690: waveform_sig_rx =-837;
15691: waveform_sig_rx =-661;
15692: waveform_sig_rx =-894;
15693: waveform_sig_rx =-948;
15694: waveform_sig_rx =-599;
15695: waveform_sig_rx =-849;
15696: waveform_sig_rx =-873;
15697: waveform_sig_rx =-743;
15698: waveform_sig_rx =-686;
15699: waveform_sig_rx =-873;
15700: waveform_sig_rx =-795;
15701: waveform_sig_rx =-630;
15702: waveform_sig_rx =-799;
15703: waveform_sig_rx =-877;
15704: waveform_sig_rx =-550;
15705: waveform_sig_rx =-698;
15706: waveform_sig_rx =-929;
15707: waveform_sig_rx =-514;
15708: waveform_sig_rx =-680;
15709: waveform_sig_rx =-854;
15710: waveform_sig_rx =-592;
15711: waveform_sig_rx =-583;
15712: waveform_sig_rx =-834;
15713: waveform_sig_rx =-603;
15714: waveform_sig_rx =-750;
15715: waveform_sig_rx =-627;
15716: waveform_sig_rx =-654;
15717: waveform_sig_rx =-673;
15718: waveform_sig_rx =-639;
15719: waveform_sig_rx =-756;
15720: waveform_sig_rx =-456;
15721: waveform_sig_rx =-822;
15722: waveform_sig_rx =-613;
15723: waveform_sig_rx =-489;
15724: waveform_sig_rx =-825;
15725: waveform_sig_rx =-583;
15726: waveform_sig_rx =-425;
15727: waveform_sig_rx =-872;
15728: waveform_sig_rx =-564;
15729: waveform_sig_rx =-377;
15730: waveform_sig_rx =-833;
15731: waveform_sig_rx =-517;
15732: waveform_sig_rx =-440;
15733: waveform_sig_rx =-672;
15734: waveform_sig_rx =-648;
15735: waveform_sig_rx =-382;
15736: waveform_sig_rx =-581;
15737: waveform_sig_rx =-589;
15738: waveform_sig_rx =-543;
15739: waveform_sig_rx =-394;
15740: waveform_sig_rx =-660;
15741: waveform_sig_rx =-568;
15742: waveform_sig_rx =-296;
15743: waveform_sig_rx =-625;
15744: waveform_sig_rx =-591;
15745: waveform_sig_rx =-263;
15746: waveform_sig_rx =-542;
15747: waveform_sig_rx =-606;
15748: waveform_sig_rx =-292;
15749: waveform_sig_rx =-465;
15750: waveform_sig_rx =-565;
15751: waveform_sig_rx =-409;
15752: waveform_sig_rx =-328;
15753: waveform_sig_rx =-554;
15754: waveform_sig_rx =-380;
15755: waveform_sig_rx =-468;
15756: waveform_sig_rx =-372;
15757: waveform_sig_rx =-445;
15758: waveform_sig_rx =-384;
15759: waveform_sig_rx =-417;
15760: waveform_sig_rx =-495;
15761: waveform_sig_rx =-152;
15762: waveform_sig_rx =-596;
15763: waveform_sig_rx =-327;
15764: waveform_sig_rx =-200;
15765: waveform_sig_rx =-629;
15766: waveform_sig_rx =-225;
15767: waveform_sig_rx =-174;
15768: waveform_sig_rx =-636;
15769: waveform_sig_rx =-191;
15770: waveform_sig_rx =-206;
15771: waveform_sig_rx =-531;
15772: waveform_sig_rx =-204;
15773: waveform_sig_rx =-237;
15774: waveform_sig_rx =-336;
15775: waveform_sig_rx =-392;
15776: waveform_sig_rx =-152;
15777: waveform_sig_rx =-258;
15778: waveform_sig_rx =-376;
15779: waveform_sig_rx =-231;
15780: waveform_sig_rx =-81;
15781: waveform_sig_rx =-450;
15782: waveform_sig_rx =-216;
15783: waveform_sig_rx =-66;
15784: waveform_sig_rx =-373;
15785: waveform_sig_rx =-245;
15786: waveform_sig_rx =-31;
15787: waveform_sig_rx =-271;
15788: waveform_sig_rx =-299;
15789: waveform_sig_rx =-55;
15790: waveform_sig_rx =-176;
15791: waveform_sig_rx =-273;
15792: waveform_sig_rx =-136;
15793: waveform_sig_rx =-11;
15794: waveform_sig_rx =-282;
15795: waveform_sig_rx =-112;
15796: waveform_sig_rx =-163;
15797: waveform_sig_rx =-107;
15798: waveform_sig_rx =-150;
15799: waveform_sig_rx =-46;
15800: waveform_sig_rx =-188;
15801: waveform_sig_rx =-157;
15802: waveform_sig_rx =118;
15803: waveform_sig_rx =-356;
15804: waveform_sig_rx =35;
15805: waveform_sig_rx =36;
15806: waveform_sig_rx =-332;
15807: waveform_sig_rx =128;
15808: waveform_sig_rx =39;
15809: waveform_sig_rx =-291;
15810: waveform_sig_rx =100;
15811: waveform_sig_rx =34;
15812: waveform_sig_rx =-169;
15813: waveform_sig_rx =29;
15814: waveform_sig_rx =64;
15815: waveform_sig_rx =-8;
15816: waveform_sig_rx =-180;
15817: waveform_sig_rx =209;
15818: waveform_sig_rx =-19;
15819: waveform_sig_rx =-138;
15820: waveform_sig_rx =130;
15821: waveform_sig_rx =125;
15822: waveform_sig_rx =-130;
15823: waveform_sig_rx =110;
15824: waveform_sig_rx =182;
15825: waveform_sig_rx =-62;
15826: waveform_sig_rx =47;
15827: waveform_sig_rx =228;
15828: waveform_sig_rx =27;
15829: waveform_sig_rx =-5;
15830: waveform_sig_rx =200;
15831: waveform_sig_rx =160;
15832: waveform_sig_rx =-11;
15833: waveform_sig_rx =130;
15834: waveform_sig_rx =335;
15835: waveform_sig_rx =-73;
15836: waveform_sig_rx =237;
15837: waveform_sig_rx =133;
15838: waveform_sig_rx =134;
15839: waveform_sig_rx =204;
15840: waveform_sig_rx =216;
15841: waveform_sig_rx =69;
15842: waveform_sig_rx =225;
15843: waveform_sig_rx =331;
15844: waveform_sig_rx =-36;
15845: waveform_sig_rx =383;
15846: waveform_sig_rx =249;
15847: waveform_sig_rx =48;
15848: waveform_sig_rx =363;
15849: waveform_sig_rx =314;
15850: waveform_sig_rx =54;
15851: waveform_sig_rx =343;
15852: waveform_sig_rx =392;
15853: waveform_sig_rx =108;
15854: waveform_sig_rx =295;
15855: waveform_sig_rx =406;
15856: waveform_sig_rx =223;
15857: waveform_sig_rx =142;
15858: waveform_sig_rx =506;
15859: waveform_sig_rx =261;
15860: waveform_sig_rx =176;
15861: waveform_sig_rx =415;
15862: waveform_sig_rx =391;
15863: waveform_sig_rx =156;
15864: waveform_sig_rx =443;
15865: waveform_sig_rx =416;
15866: waveform_sig_rx =262;
15867: waveform_sig_rx =317;
15868: waveform_sig_rx =468;
15869: waveform_sig_rx =390;
15870: waveform_sig_rx =209;
15871: waveform_sig_rx =547;
15872: waveform_sig_rx =459;
15873: waveform_sig_rx =185;
15874: waveform_sig_rx =521;
15875: waveform_sig_rx =533;
15876: waveform_sig_rx =211;
15877: waveform_sig_rx =596;
15878: waveform_sig_rx =337;
15879: waveform_sig_rx =486;
15880: waveform_sig_rx =473;
15881: waveform_sig_rx =462;
15882: waveform_sig_rx =391;
15883: waveform_sig_rx =473;
15884: waveform_sig_rx =577;
15885: waveform_sig_rx =284;
15886: waveform_sig_rx =617;
15887: waveform_sig_rx =531;
15888: waveform_sig_rx =310;
15889: waveform_sig_rx =614;
15890: waveform_sig_rx =603;
15891: waveform_sig_rx =300;
15892: waveform_sig_rx =596;
15893: waveform_sig_rx =648;
15894: waveform_sig_rx =350;
15895: waveform_sig_rx =567;
15896: waveform_sig_rx =699;
15897: waveform_sig_rx =441;
15898: waveform_sig_rx =453;
15899: waveform_sig_rx =791;
15900: waveform_sig_rx =457;
15901: waveform_sig_rx =500;
15902: waveform_sig_rx =676;
15903: waveform_sig_rx =635;
15904: waveform_sig_rx =489;
15905: waveform_sig_rx =646;
15906: waveform_sig_rx =707;
15907: waveform_sig_rx =532;
15908: waveform_sig_rx =529;
15909: waveform_sig_rx =816;
15910: waveform_sig_rx =600;
15911: waveform_sig_rx =471;
15912: waveform_sig_rx =854;
15913: waveform_sig_rx =631;
15914: waveform_sig_rx =489;
15915: waveform_sig_rx =817;
15916: waveform_sig_rx =709;
15917: waveform_sig_rx =535;
15918: waveform_sig_rx =787;
15919: waveform_sig_rx =556;
15920: waveform_sig_rx =796;
15921: waveform_sig_rx =645;
15922: waveform_sig_rx =763;
15923: waveform_sig_rx =659;
15924: waveform_sig_rx =710;
15925: waveform_sig_rx =861;
15926: waveform_sig_rx =526;
15927: waveform_sig_rx =850;
15928: waveform_sig_rx =798;
15929: waveform_sig_rx =553;
15930: waveform_sig_rx =870;
15931: waveform_sig_rx =845;
15932: waveform_sig_rx =525;
15933: waveform_sig_rx =840;
15934: waveform_sig_rx =924;
15935: waveform_sig_rx =523;
15936: waveform_sig_rx =859;
15937: waveform_sig_rx =931;
15938: waveform_sig_rx =596;
15939: waveform_sig_rx =788;
15940: waveform_sig_rx =950;
15941: waveform_sig_rx =707;
15942: waveform_sig_rx =780;
15943: waveform_sig_rx =819;
15944: waveform_sig_rx =943;
15945: waveform_sig_rx =625;
15946: waveform_sig_rx =861;
15947: waveform_sig_rx =983;
15948: waveform_sig_rx =667;
15949: waveform_sig_rx =826;
15950: waveform_sig_rx =1028;
15951: waveform_sig_rx =762;
15952: waveform_sig_rx =741;
15953: waveform_sig_rx =1058;
15954: waveform_sig_rx =846;
15955: waveform_sig_rx =713;
15956: waveform_sig_rx =1022;
15957: waveform_sig_rx =910;
15958: waveform_sig_rx =767;
15959: waveform_sig_rx =997;
15960: waveform_sig_rx =762;
15961: waveform_sig_rx =1037;
15962: waveform_sig_rx =807;
15963: waveform_sig_rx =1012;
15964: waveform_sig_rx =853;
15965: waveform_sig_rx =892;
15966: waveform_sig_rx =1083;
15967: waveform_sig_rx =685;
15968: waveform_sig_rx =1071;
15969: waveform_sig_rx =1035;
15970: waveform_sig_rx =692;
15971: waveform_sig_rx =1138;
15972: waveform_sig_rx =1020;
15973: waveform_sig_rx =684;
15974: waveform_sig_rx =1155;
15975: waveform_sig_rx =1022;
15976: waveform_sig_rx =752;
15977: waveform_sig_rx =1108;
15978: waveform_sig_rx =1036;
15979: waveform_sig_rx =857;
15980: waveform_sig_rx =959;
15981: waveform_sig_rx =1107;
15982: waveform_sig_rx =939;
15983: waveform_sig_rx =899;
15984: waveform_sig_rx =1047;
15985: waveform_sig_rx =1118;
15986: waveform_sig_rx =788;
15987: waveform_sig_rx =1111;
15988: waveform_sig_rx =1114;
15989: waveform_sig_rx =830;
15990: waveform_sig_rx =1028;
15991: waveform_sig_rx =1182;
15992: waveform_sig_rx =916;
15993: waveform_sig_rx =938;
15994: waveform_sig_rx =1198;
15995: waveform_sig_rx =976;
15996: waveform_sig_rx =906;
15997: waveform_sig_rx =1144;
15998: waveform_sig_rx =1075;
15999: waveform_sig_rx =941;
16000: waveform_sig_rx =1089;
16001: waveform_sig_rx =973;
16002: waveform_sig_rx =1158;
16003: waveform_sig_rx =942;
16004: waveform_sig_rx =1205;
16005: waveform_sig_rx =887;
16006: waveform_sig_rx =1106;
16007: waveform_sig_rx =1213;
16008: waveform_sig_rx =777;
16009: waveform_sig_rx =1298;
16010: waveform_sig_rx =1056;
16011: waveform_sig_rx =835;
16012: waveform_sig_rx =1309;
16013: waveform_sig_rx =1057;
16014: waveform_sig_rx =884;
16015: waveform_sig_rx =1240;
16016: waveform_sig_rx =1124;
16017: waveform_sig_rx =909;
16018: waveform_sig_rx =1185;
16019: waveform_sig_rx =1176;
16020: waveform_sig_rx =969;
16021: waveform_sig_rx =1035;
16022: waveform_sig_rx =1251;
16023: waveform_sig_rx =1045;
16024: waveform_sig_rx =996;
16025: waveform_sig_rx =1204;
16026: waveform_sig_rx =1198;
16027: waveform_sig_rx =873;
16028: waveform_sig_rx =1261;
16029: waveform_sig_rx =1185;
16030: waveform_sig_rx =933;
16031: waveform_sig_rx =1163;
16032: waveform_sig_rx =1219;
16033: waveform_sig_rx =1026;
16034: waveform_sig_rx =1054;
16035: waveform_sig_rx =1250;
16036: waveform_sig_rx =1106;
16037: waveform_sig_rx =982;
16038: waveform_sig_rx =1239;
16039: waveform_sig_rx =1208;
16040: waveform_sig_rx =942;
16041: waveform_sig_rx =1239;
16042: waveform_sig_rx =1067;
16043: waveform_sig_rx =1167;
16044: waveform_sig_rx =1104;
16045: waveform_sig_rx =1246;
16046: waveform_sig_rx =966;
16047: waveform_sig_rx =1268;
16048: waveform_sig_rx =1194;
16049: waveform_sig_rx =902;
16050: waveform_sig_rx =1378;
16051: waveform_sig_rx =1069;
16052: waveform_sig_rx =1007;
16053: waveform_sig_rx =1323;
16054: waveform_sig_rx =1147;
16055: waveform_sig_rx =957;
16056: waveform_sig_rx =1281;
16057: waveform_sig_rx =1184;
16058: waveform_sig_rx =956;
16059: waveform_sig_rx =1223;
16060: waveform_sig_rx =1228;
16061: waveform_sig_rx =1027;
16062: waveform_sig_rx =1098;
16063: waveform_sig_rx =1317;
16064: waveform_sig_rx =1075;
16065: waveform_sig_rx =1034;
16066: waveform_sig_rx =1287;
16067: waveform_sig_rx =1177;
16068: waveform_sig_rx =936;
16069: waveform_sig_rx =1309;
16070: waveform_sig_rx =1129;
16071: waveform_sig_rx =1051;
16072: waveform_sig_rx =1160;
16073: waveform_sig_rx =1249;
16074: waveform_sig_rx =1122;
16075: waveform_sig_rx =999;
16076: waveform_sig_rx =1342;
16077: waveform_sig_rx =1123;
16078: waveform_sig_rx =961;
16079: waveform_sig_rx =1340;
16080: waveform_sig_rx =1151;
16081: waveform_sig_rx =1001;
16082: waveform_sig_rx =1301;
16083: waveform_sig_rx =1018;
16084: waveform_sig_rx =1245;
16085: waveform_sig_rx =1094;
16086: waveform_sig_rx =1206;
16087: waveform_sig_rx =992;
16088: waveform_sig_rx =1248;
16089: waveform_sig_rx =1171;
16090: waveform_sig_rx =960;
16091: waveform_sig_rx =1335;
16092: waveform_sig_rx =1072;
16093: waveform_sig_rx =1001;
16094: waveform_sig_rx =1297;
16095: waveform_sig_rx =1115;
16096: waveform_sig_rx =948;
16097: waveform_sig_rx =1235;
16098: waveform_sig_rx =1192;
16099: waveform_sig_rx =942;
16100: waveform_sig_rx =1192;
16101: waveform_sig_rx =1255;
16102: waveform_sig_rx =938;
16103: waveform_sig_rx =1127;
16104: waveform_sig_rx =1300;
16105: waveform_sig_rx =980;
16106: waveform_sig_rx =1092;
16107: waveform_sig_rx =1231;
16108: waveform_sig_rx =1123;
16109: waveform_sig_rx =985;
16110: waveform_sig_rx =1224;
16111: waveform_sig_rx =1160;
16112: waveform_sig_rx =996;
16113: waveform_sig_rx =1067;
16114: waveform_sig_rx =1263;
16115: waveform_sig_rx =1000;
16116: waveform_sig_rx =979;
16117: waveform_sig_rx =1320;
16118: waveform_sig_rx =983;
16119: waveform_sig_rx =937;
16120: waveform_sig_rx =1278;
16121: waveform_sig_rx =1051;
16122: waveform_sig_rx =988;
16123: waveform_sig_rx =1197;
16124: waveform_sig_rx =930;
16125: waveform_sig_rx =1207;
16126: waveform_sig_rx =988;
16127: waveform_sig_rx =1146;
16128: waveform_sig_rx =941;
16129: waveform_sig_rx =1141;
16130: waveform_sig_rx =1105;
16131: waveform_sig_rx =873;
16132: waveform_sig_rx =1217;
16133: waveform_sig_rx =1023;
16134: waveform_sig_rx =887;
16135: waveform_sig_rx =1221;
16136: waveform_sig_rx =1050;
16137: waveform_sig_rx =838;
16138: waveform_sig_rx =1223;
16139: waveform_sig_rx =1072;
16140: waveform_sig_rx =827;
16141: waveform_sig_rx =1138;
16142: waveform_sig_rx =1122;
16143: waveform_sig_rx =811;
16144: waveform_sig_rx =1060;
16145: waveform_sig_rx =1136;
16146: waveform_sig_rx =869;
16147: waveform_sig_rx =987;
16148: waveform_sig_rx =1061;
16149: waveform_sig_rx =1031;
16150: waveform_sig_rx =843;
16151: waveform_sig_rx =1078;
16152: waveform_sig_rx =1068;
16153: waveform_sig_rx =823;
16154: waveform_sig_rx =995;
16155: waveform_sig_rx =1159;
16156: waveform_sig_rx =802;
16157: waveform_sig_rx =930;
16158: waveform_sig_rx =1165;
16159: waveform_sig_rx =826;
16160: waveform_sig_rx =892;
16161: waveform_sig_rx =1096;
16162: waveform_sig_rx =922;
16163: waveform_sig_rx =872;
16164: waveform_sig_rx =1003;
16165: waveform_sig_rx =842;
16166: waveform_sig_rx =1068;
16167: waveform_sig_rx =809;
16168: waveform_sig_rx =1046;
16169: waveform_sig_rx =767;
16170: waveform_sig_rx =996;
16171: waveform_sig_rx =981;
16172: waveform_sig_rx =679;
16173: waveform_sig_rx =1085;
16174: waveform_sig_rx =884;
16175: waveform_sig_rx =695;
16176: waveform_sig_rx =1112;
16177: waveform_sig_rx =853;
16178: waveform_sig_rx =636;
16179: waveform_sig_rx =1119;
16180: waveform_sig_rx =842;
16181: waveform_sig_rx =706;
16182: waveform_sig_rx =1001;
16183: waveform_sig_rx =886;
16184: waveform_sig_rx =696;
16185: waveform_sig_rx =874;
16186: waveform_sig_rx =935;
16187: waveform_sig_rx =742;
16188: waveform_sig_rx =789;
16189: waveform_sig_rx =915;
16190: waveform_sig_rx =878;
16191: waveform_sig_rx =627;
16192: waveform_sig_rx =946;
16193: waveform_sig_rx =900;
16194: waveform_sig_rx =592;
16195: waveform_sig_rx =897;
16196: waveform_sig_rx =918;
16197: waveform_sig_rx =588;
16198: waveform_sig_rx =801;
16199: waveform_sig_rx =900;
16200: waveform_sig_rx =678;
16201: waveform_sig_rx =683;
16202: waveform_sig_rx =857;
16203: waveform_sig_rx =791;
16204: waveform_sig_rx =642;
16205: waveform_sig_rx =828;
16206: waveform_sig_rx =658;
16207: waveform_sig_rx =813;
16208: waveform_sig_rx =659;
16209: waveform_sig_rx =847;
16210: waveform_sig_rx =533;
16211: waveform_sig_rx =847;
16212: waveform_sig_rx =713;
16213: waveform_sig_rx =487;
16214: waveform_sig_rx =903;
16215: waveform_sig_rx =609;
16216: waveform_sig_rx =482;
16217: waveform_sig_rx =926;
16218: waveform_sig_rx =582;
16219: waveform_sig_rx =465;
16220: waveform_sig_rx =921;
16221: waveform_sig_rx =521;
16222: waveform_sig_rx =570;
16223: waveform_sig_rx =742;
16224: waveform_sig_rx =650;
16225: waveform_sig_rx =532;
16226: waveform_sig_rx =577;
16227: waveform_sig_rx =765;
16228: waveform_sig_rx =510;
16229: waveform_sig_rx =492;
16230: waveform_sig_rx =778;
16231: waveform_sig_rx =581;
16232: waveform_sig_rx =415;
16233: waveform_sig_rx =794;
16234: waveform_sig_rx =578;
16235: waveform_sig_rx =423;
16236: waveform_sig_rx =624;
16237: waveform_sig_rx =620;
16238: waveform_sig_rx =394;
16239: waveform_sig_rx =507;
16240: waveform_sig_rx =653;
16241: waveform_sig_rx =430;
16242: waveform_sig_rx =395;
16243: waveform_sig_rx =654;
16244: waveform_sig_rx =502;
16245: waveform_sig_rx =365;
16246: waveform_sig_rx =573;
16247: waveform_sig_rx =377;
16248: waveform_sig_rx =524;
16249: waveform_sig_rx =412;
16250: waveform_sig_rx =541;
16251: waveform_sig_rx =255;
16252: waveform_sig_rx =627;
16253: waveform_sig_rx =391;
16254: waveform_sig_rx =254;
16255: waveform_sig_rx =693;
16256: waveform_sig_rx =263;
16257: waveform_sig_rx =304;
16258: waveform_sig_rx =678;
16259: waveform_sig_rx =255;
16260: waveform_sig_rx =301;
16261: waveform_sig_rx =560;
16262: waveform_sig_rx =289;
16263: waveform_sig_rx =315;
16264: waveform_sig_rx =404;
16265: waveform_sig_rx =465;
16266: waveform_sig_rx =170;
16267: waveform_sig_rx =333;
16268: waveform_sig_rx =531;
16269: waveform_sig_rx =141;
16270: waveform_sig_rx =294;
16271: waveform_sig_rx =453;
16272: waveform_sig_rx =228;
16273: waveform_sig_rx =198;
16274: waveform_sig_rx =413;
16275: waveform_sig_rx =292;
16276: waveform_sig_rx =141;
16277: waveform_sig_rx =327;
16278: waveform_sig_rx =364;
16279: waveform_sig_rx =99;
16280: waveform_sig_rx =221;
16281: waveform_sig_rx =372;
16282: waveform_sig_rx =142;
16283: waveform_sig_rx =107;
16284: waveform_sig_rx =397;
16285: waveform_sig_rx =192;
16286: waveform_sig_rx =76;
16287: waveform_sig_rx =317;
16288: waveform_sig_rx =58;
16289: waveform_sig_rx =257;
16290: waveform_sig_rx =145;
16291: waveform_sig_rx =208;
16292: waveform_sig_rx =-15;
16293: waveform_sig_rx =348;
16294: waveform_sig_rx =45;
16295: waveform_sig_rx =28;
16296: waveform_sig_rx =336;
16297: waveform_sig_rx =-23;
16298: waveform_sig_rx =58;
16299: waveform_sig_rx =273;
16300: waveform_sig_rx =27;
16301: waveform_sig_rx =-48;
16302: waveform_sig_rx =264;
16303: waveform_sig_rx =37;
16304: waveform_sig_rx =-101;
16305: waveform_sig_rx =165;
16306: waveform_sig_rx =130;
16307: waveform_sig_rx =-201;
16308: waveform_sig_rx =134;
16309: waveform_sig_rx =149;
16310: waveform_sig_rx =-134;
16311: waveform_sig_rx =38;
16312: waveform_sig_rx =105;
16313: waveform_sig_rx =-21;
16314: waveform_sig_rx =-120;
16315: waveform_sig_rx =124;
16316: waveform_sig_rx =6;
16317: waveform_sig_rx =-163;
16318: waveform_sig_rx =31;
16319: waveform_sig_rx =75;
16320: waveform_sig_rx =-207;
16321: waveform_sig_rx =-112;
16322: waveform_sig_rx =110;
16323: waveform_sig_rx =-195;
16324: waveform_sig_rx =-206;
16325: waveform_sig_rx =137;
16326: waveform_sig_rx =-220;
16327: waveform_sig_rx =-146;
16328: waveform_sig_rx =-11;
16329: waveform_sig_rx =-287;
16330: waveform_sig_rx =37;
16331: waveform_sig_rx =-232;
16332: waveform_sig_rx =-70;
16333: waveform_sig_rx =-256;
16334: waveform_sig_rx =-23;
16335: waveform_sig_rx =-213;
16336: waveform_sig_rx =-286;
16337: waveform_sig_rx =-18;
16338: waveform_sig_rx =-264;
16339: waveform_sig_rx =-327;
16340: waveform_sig_rx =16;
16341: waveform_sig_rx =-308;
16342: waveform_sig_rx =-402;
16343: waveform_sig_rx =22;
16344: waveform_sig_rx =-328;
16345: waveform_sig_rx =-365;
16346: waveform_sig_rx =-114;
16347: waveform_sig_rx =-234;
16348: waveform_sig_rx =-467;
16349: waveform_sig_rx =-165;
16350: waveform_sig_rx =-196;
16351: waveform_sig_rx =-407;
16352: waveform_sig_rx =-284;
16353: waveform_sig_rx =-203;
16354: waveform_sig_rx =-340;
16355: waveform_sig_rx =-426;
16356: waveform_sig_rx =-209;
16357: waveform_sig_rx =-292;
16358: waveform_sig_rx =-488;
16359: waveform_sig_rx =-277;
16360: waveform_sig_rx =-194;
16361: waveform_sig_rx =-578;
16362: waveform_sig_rx =-313;
16363: waveform_sig_rx =-202;
16364: waveform_sig_rx =-564;
16365: waveform_sig_rx =-400;
16366: waveform_sig_rx =-248;
16367: waveform_sig_rx =-493;
16368: waveform_sig_rx =-409;
16369: waveform_sig_rx =-410;
16370: waveform_sig_rx =-473;
16371: waveform_sig_rx =-318;
16372: waveform_sig_rx =-541;
16373: waveform_sig_rx =-311;
16374: waveform_sig_rx =-623;
16375: waveform_sig_rx =-294;
16376: waveform_sig_rx =-516;
16377: waveform_sig_rx =-624;
16378: waveform_sig_rx =-252;
16379: waveform_sig_rx =-609;
16380: waveform_sig_rx =-631;
16381: waveform_sig_rx =-247;
16382: waveform_sig_rx =-637;
16383: waveform_sig_rx =-659;
16384: waveform_sig_rx =-268;
16385: waveform_sig_rx =-651;
16386: waveform_sig_rx =-653;
16387: waveform_sig_rx =-373;
16388: waveform_sig_rx =-556;
16389: waveform_sig_rx =-740;
16390: waveform_sig_rx =-451;
16391: waveform_sig_rx =-525;
16392: waveform_sig_rx =-673;
16393: waveform_sig_rx =-633;
16394: waveform_sig_rx =-474;
16395: waveform_sig_rx =-611;
16396: waveform_sig_rx =-768;
16397: waveform_sig_rx =-433;
16398: waveform_sig_rx =-604;
16399: waveform_sig_rx =-812;
16400: waveform_sig_rx =-484;
16401: waveform_sig_rx =-545;
16402: waveform_sig_rx =-830;
16403: waveform_sig_rx =-575;
16404: waveform_sig_rx =-546;
16405: waveform_sig_rx =-769;
16406: waveform_sig_rx =-679;
16407: waveform_sig_rx =-544;
16408: waveform_sig_rx =-712;
16409: waveform_sig_rx =-740;
16410: waveform_sig_rx =-677;
16411: waveform_sig_rx =-701;
16412: waveform_sig_rx =-666;
16413: waveform_sig_rx =-756;
16414: waveform_sig_rx =-613;
16415: waveform_sig_rx =-936;
16416: waveform_sig_rx =-483;
16417: waveform_sig_rx =-842;
16418: waveform_sig_rx =-865;
16419: waveform_sig_rx =-489;
16420: waveform_sig_rx =-909;
16421: waveform_sig_rx =-830;
16422: waveform_sig_rx =-516;
16423: waveform_sig_rx =-936;
16424: waveform_sig_rx =-875;
16425: waveform_sig_rx =-526;
16426: waveform_sig_rx =-937;
16427: waveform_sig_rx =-848;
16428: waveform_sig_rx =-663;
16429: waveform_sig_rx =-821;
16430: waveform_sig_rx =-926;
16431: waveform_sig_rx =-745;
16432: waveform_sig_rx =-728;
16433: waveform_sig_rx =-902;
16434: waveform_sig_rx =-921;
16435: waveform_sig_rx =-644;
16436: waveform_sig_rx =-925;
16437: waveform_sig_rx =-985;
16438: waveform_sig_rx =-622;
16439: waveform_sig_rx =-940;
16440: waveform_sig_rx =-993;
16441: waveform_sig_rx =-733;
16442: waveform_sig_rx =-822;
16443: waveform_sig_rx =-1014;
16444: waveform_sig_rx =-830;
16445: waveform_sig_rx =-762;
16446: waveform_sig_rx =-1006;
16447: waveform_sig_rx =-942;
16448: waveform_sig_rx =-747;
16449: waveform_sig_rx =-954;
16450: waveform_sig_rx =-952;
16451: waveform_sig_rx =-865;
16452: waveform_sig_rx =-935;
16453: waveform_sig_rx =-892;
16454: waveform_sig_rx =-933;
16455: waveform_sig_rx =-877;
16456: waveform_sig_rx =-1136;
16457: waveform_sig_rx =-680;
16458: waveform_sig_rx =-1114;
16459: waveform_sig_rx =-1006;
16460: waveform_sig_rx =-709;
16461: waveform_sig_rx =-1194;
16462: waveform_sig_rx =-947;
16463: waveform_sig_rx =-776;
16464: waveform_sig_rx =-1138;
16465: waveform_sig_rx =-1029;
16466: waveform_sig_rx =-799;
16467: waveform_sig_rx =-1092;
16468: waveform_sig_rx =-1069;
16469: waveform_sig_rx =-870;
16470: waveform_sig_rx =-976;
16471: waveform_sig_rx =-1175;
16472: waveform_sig_rx =-904;
16473: waveform_sig_rx =-920;
16474: waveform_sig_rx =-1120;
16475: waveform_sig_rx =-1062;
16476: waveform_sig_rx =-825;
16477: waveform_sig_rx =-1149;
16478: waveform_sig_rx =-1121;
16479: waveform_sig_rx =-821;
16480: waveform_sig_rx =-1145;
16481: waveform_sig_rx =-1117;
16482: waveform_sig_rx =-958;
16483: waveform_sig_rx =-1004;
16484: waveform_sig_rx =-1173;
16485: waveform_sig_rx =-1053;
16486: waveform_sig_rx =-892;
16487: waveform_sig_rx =-1192;
16488: waveform_sig_rx =-1129;
16489: waveform_sig_rx =-835;
16490: waveform_sig_rx =-1209;
16491: waveform_sig_rx =-1095;
16492: waveform_sig_rx =-1019;
16493: waveform_sig_rx =-1145;
16494: waveform_sig_rx =-1014;
16495: waveform_sig_rx =-1086;
16496: waveform_sig_rx =-1065;
16497: waveform_sig_rx =-1227;
16498: waveform_sig_rx =-850;
16499: waveform_sig_rx =-1300;
16500: waveform_sig_rx =-1088;
16501: waveform_sig_rx =-935;
16502: waveform_sig_rx =-1289;
16503: waveform_sig_rx =-1083;
16504: waveform_sig_rx =-957;
16505: waveform_sig_rx =-1230;
16506: waveform_sig_rx =-1181;
16507: waveform_sig_rx =-928;
16508: waveform_sig_rx =-1198;
16509: waveform_sig_rx =-1204;
16510: waveform_sig_rx =-993;
16511: waveform_sig_rx =-1096;
16512: waveform_sig_rx =-1337;
16513: waveform_sig_rx =-988;
16514: waveform_sig_rx =-1046;
16515: waveform_sig_rx =-1274;
16516: waveform_sig_rx =-1128;
16517: waveform_sig_rx =-990;
16518: waveform_sig_rx =-1290;
16519: waveform_sig_rx =-1161;
16520: waveform_sig_rx =-1016;
16521: waveform_sig_rx =-1212;
16522: waveform_sig_rx =-1203;
16523: waveform_sig_rx =-1086;
16524: waveform_sig_rx =-1046;
16525: waveform_sig_rx =-1324;
16526: waveform_sig_rx =-1131;
16527: waveform_sig_rx =-966;
16528: waveform_sig_rx =-1352;
16529: waveform_sig_rx =-1149;
16530: waveform_sig_rx =-955;
16531: waveform_sig_rx =-1329;
16532: waveform_sig_rx =-1113;
16533: waveform_sig_rx =-1165;
16534: waveform_sig_rx =-1224;
16535: waveform_sig_rx =-1084;
16536: waveform_sig_rx =-1213;
16537: waveform_sig_rx =-1134;
16538: waveform_sig_rx =-1277;
16539: waveform_sig_rx =-955;
16540: waveform_sig_rx =-1327;
16541: waveform_sig_rx =-1148;
16542: waveform_sig_rx =-1012;
16543: waveform_sig_rx =-1332;
16544: waveform_sig_rx =-1162;
16545: waveform_sig_rx =-1017;
16546: waveform_sig_rx =-1288;
16547: waveform_sig_rx =-1254;
16548: waveform_sig_rx =-948;
16549: waveform_sig_rx =-1293;
16550: waveform_sig_rx =-1268;
16551: waveform_sig_rx =-984;
16552: waveform_sig_rx =-1198;
16553: waveform_sig_rx =-1366;
16554: waveform_sig_rx =-991;
16555: waveform_sig_rx =-1164;
16556: waveform_sig_rx =-1284;
16557: waveform_sig_rx =-1145;
16558: waveform_sig_rx =-1069;
16559: waveform_sig_rx =-1259;
16560: waveform_sig_rx =-1205;
16561: waveform_sig_rx =-1042;
16562: waveform_sig_rx =-1196;
16563: waveform_sig_rx =-1304;
16564: waveform_sig_rx =-1047;
16565: waveform_sig_rx =-1068;
16566: waveform_sig_rx =-1391;
16567: waveform_sig_rx =-1056;
16568: waveform_sig_rx =-1051;
16569: waveform_sig_rx =-1344;
16570: waveform_sig_rx =-1109;
16571: waveform_sig_rx =-1007;
16572: waveform_sig_rx =-1297;
16573: waveform_sig_rx =-1092;
16574: waveform_sig_rx =-1184;
16575: waveform_sig_rx =-1177;
16576: waveform_sig_rx =-1087;
16577: waveform_sig_rx =-1202;
16578: waveform_sig_rx =-1102;
16579: waveform_sig_rx =-1263;
16580: waveform_sig_rx =-971;
16581: waveform_sig_rx =-1282;
16582: waveform_sig_rx =-1167;
16583: waveform_sig_rx =-994;
16584: waveform_sig_rx =-1279;
16585: waveform_sig_rx =-1175;
16586: waveform_sig_rx =-924;
16587: waveform_sig_rx =-1291;
16588: waveform_sig_rx =-1206;
16589: waveform_sig_rx =-831;
16590: waveform_sig_rx =-1318;
16591: waveform_sig_rx =-1154;
16592: waveform_sig_rx =-940;
16593: waveform_sig_rx =-1207;
16594: waveform_sig_rx =-1249;
16595: waveform_sig_rx =-959;
16596: waveform_sig_rx =-1152;
16597: waveform_sig_rx =-1175;
16598: waveform_sig_rx =-1125;
16599: waveform_sig_rx =-992;
16600: waveform_sig_rx =-1204;
16601: waveform_sig_rx =-1213;
16602: waveform_sig_rx =-921;
16603: waveform_sig_rx =-1143;
16604: waveform_sig_rx =-1254;
16605: waveform_sig_rx =-935;
16606: waveform_sig_rx =-1045;
16607: waveform_sig_rx =-1306;
16608: waveform_sig_rx =-941;
16609: waveform_sig_rx =-1023;
16610: waveform_sig_rx =-1238;
16611: waveform_sig_rx =-1025;
16612: waveform_sig_rx =-982;
16613: waveform_sig_rx =-1179;
16614: waveform_sig_rx =-1026;
16615: waveform_sig_rx =-1115;
16616: waveform_sig_rx =-1017;
16617: waveform_sig_rx =-1063;
16618: waveform_sig_rx =-1083;
16619: waveform_sig_rx =-994;
16620: waveform_sig_rx =-1223;
16621: waveform_sig_rx =-813;
16622: waveform_sig_rx =-1206;
16623: waveform_sig_rx =-1076;
16624: waveform_sig_rx =-812;
16625: waveform_sig_rx =-1243;
16626: waveform_sig_rx =-1014;
16627: waveform_sig_rx =-787;
16628: waveform_sig_rx =-1265;
16629: waveform_sig_rx =-1014;
16630: waveform_sig_rx =-791;
16631: waveform_sig_rx =-1228;
16632: waveform_sig_rx =-989;
16633: waveform_sig_rx =-886;
16634: waveform_sig_rx =-1071;
16635: waveform_sig_rx =-1113;
16636: waveform_sig_rx =-842;
16637: waveform_sig_rx =-981;
16638: waveform_sig_rx =-1049;
16639: waveform_sig_rx =-1003;
16640: waveform_sig_rx =-808;
16641: waveform_sig_rx =-1090;
16642: waveform_sig_rx =-1047;
16643: waveform_sig_rx =-760;
16644: waveform_sig_rx =-1090;
16645: waveform_sig_rx =-1068;
16646: waveform_sig_rx =-768;
16647: waveform_sig_rx =-999;
16648: waveform_sig_rx =-1089;
16649: waveform_sig_rx =-838;
16650: waveform_sig_rx =-909;
16651: waveform_sig_rx =-1025;
16652: waveform_sig_rx =-958;
16653: waveform_sig_rx =-758;
16654: waveform_sig_rx =-1023;
16655: waveform_sig_rx =-917;
16656: waveform_sig_rx =-898;
16657: waveform_sig_rx =-900;
16658: waveform_sig_rx =-901;
16659: waveform_sig_rx =-854;
16660: waveform_sig_rx =-876;
16661: waveform_sig_rx =-1021;
16662: waveform_sig_rx =-617;
16663: waveform_sig_rx =-1114;
16664: waveform_sig_rx =-835;
16665: waveform_sig_rx =-663;
16666: waveform_sig_rx =-1113;
16667: waveform_sig_rx =-768;
16668: waveform_sig_rx =-664;
16669: waveform_sig_rx =-1093;
16670: waveform_sig_rx =-765;
16671: waveform_sig_rx =-686;
16672: waveform_sig_rx =-1011;
16673: waveform_sig_rx =-786;
16674: waveform_sig_rx =-735;
16675: waveform_sig_rx =-841;
16676: waveform_sig_rx =-960;
16677: waveform_sig_rx =-682;
16678: waveform_sig_rx =-757;
16679: waveform_sig_rx =-926;
16680: waveform_sig_rx =-783;
16681: waveform_sig_rx =-614;
16682: waveform_sig_rx =-965;
16683: waveform_sig_rx =-795;
16684: waveform_sig_rx =-579;
16685: waveform_sig_rx =-908;
16686: waveform_sig_rx =-800;
16687: waveform_sig_rx =-615;
16688: waveform_sig_rx =-781;
16689: waveform_sig_rx =-838;
16690: waveform_sig_rx =-670;
16691: waveform_sig_rx =-631;
16692: waveform_sig_rx =-847;
16693: waveform_sig_rx =-750;
16694: waveform_sig_rx =-504;
16695: waveform_sig_rx =-886;
16696: waveform_sig_rx =-646;
16697: waveform_sig_rx =-680;
16698: waveform_sig_rx =-729;
16699: waveform_sig_rx =-647;
16700: waveform_sig_rx =-653;
16701: waveform_sig_rx =-702;
16702: waveform_sig_rx =-749;
16703: waveform_sig_rx =-436;
16704: waveform_sig_rx =-897;
16705: waveform_sig_rx =-555;
16706: waveform_sig_rx =-485;
16707: waveform_sig_rx =-880;
16708: waveform_sig_rx =-493;
16709: waveform_sig_rx =-502;
16710: waveform_sig_rx =-825;
16711: waveform_sig_rx =-517;
16712: waveform_sig_rx =-500;
16713: waveform_sig_rx =-700;
16714: waveform_sig_rx =-587;
16715: waveform_sig_rx =-482;
16716: waveform_sig_rx =-529;
16717: waveform_sig_rx =-788;
16718: waveform_sig_rx =-353;
16719: waveform_sig_rx =-560;
16720: waveform_sig_rx =-706;
16721: waveform_sig_rx =-441;
16722: waveform_sig_rx =-460;
16723: waveform_sig_rx =-687;
16724: waveform_sig_rx =-503;
16725: waveform_sig_rx =-408;
16726: waveform_sig_rx =-597;
16727: waveform_sig_rx =-581;
16728: waveform_sig_rx =-369;
16729: waveform_sig_rx =-492;
16730: waveform_sig_rx =-653;
16731: waveform_sig_rx =-376;
16732: waveform_sig_rx =-401;
16733: waveform_sig_rx =-614;
16734: waveform_sig_rx =-447;
16735: waveform_sig_rx =-250;
16736: waveform_sig_rx =-647;
16737: waveform_sig_rx =-351;
16738: waveform_sig_rx =-423;
16739: waveform_sig_rx =-476;
16740: waveform_sig_rx =-332;
16741: waveform_sig_rx =-398;
16742: waveform_sig_rx =-453;
16743: waveform_sig_rx =-410;
16744: waveform_sig_rx =-224;
16745: waveform_sig_rx =-599;
16746: waveform_sig_rx =-265;
16747: waveform_sig_rx =-305;
16748: waveform_sig_rx =-518;
16749: waveform_sig_rx =-280;
16750: waveform_sig_rx =-236;
16751: waveform_sig_rx =-499;
16752: waveform_sig_rx =-331;
16753: waveform_sig_rx =-139;
16754: waveform_sig_rx =-470;
16755: waveform_sig_rx =-351;
16756: waveform_sig_rx =-142;
16757: waveform_sig_rx =-370;
16758: waveform_sig_rx =-450;
16759: waveform_sig_rx =-48;
16760: waveform_sig_rx =-361;
16761: waveform_sig_rx =-362;
16762: waveform_sig_rx =-200;
16763: waveform_sig_rx =-187;
16764: waveform_sig_rx =-358;
16765: waveform_sig_rx =-241;
16766: waveform_sig_rx =-103;
16767: waveform_sig_rx =-303;
16768: waveform_sig_rx =-332;
16769: waveform_sig_rx =-54;
16770: waveform_sig_rx =-186;
16771: waveform_sig_rx =-368;
16772: waveform_sig_rx =-48;
16773: waveform_sig_rx =-95;
16774: waveform_sig_rx =-369;
16775: waveform_sig_rx =-87;
16776: waveform_sig_rx =-4;
16777: waveform_sig_rx =-378;
16778: waveform_sig_rx =-1;
16779: waveform_sig_rx =-226;
16780: waveform_sig_rx =-122;
16781: waveform_sig_rx =-66;
16782: waveform_sig_rx =-169;
16783: waveform_sig_rx =-105;
16784: waveform_sig_rx =-167;
16785: waveform_sig_rx =46;
16786: waveform_sig_rx =-241;
16787: waveform_sig_rx =-37;
16788: waveform_sig_rx =59;
16789: waveform_sig_rx =-260;
16790: waveform_sig_rx =-14;
16791: waveform_sig_rx =141;
16792: waveform_sig_rx =-296;
16793: waveform_sig_rx =24;
16794: waveform_sig_rx =162;
16795: waveform_sig_rx =-249;
16796: waveform_sig_rx =29;
16797: waveform_sig_rx =136;
16798: waveform_sig_rx =-104;
16799: waveform_sig_rx =-113;
16800: waveform_sig_rx =197;
16801: waveform_sig_rx =-50;
16802: waveform_sig_rx =-61;
16803: waveform_sig_rx =61;
16804: waveform_sig_rx =142;
16805: waveform_sig_rx =-75;
16806: waveform_sig_rx =46;
16807: waveform_sig_rx =219;
16808: waveform_sig_rx =-17;
16809: waveform_sig_rx =-52;
16810: waveform_sig_rx =291;
16811: waveform_sig_rx =76;
16812: waveform_sig_rx =-110;
16813: waveform_sig_rx =322;
16814: waveform_sig_rx =126;
16815: waveform_sig_rx =-25;
16816: waveform_sig_rx =264;
16817: waveform_sig_rx =188;
16818: waveform_sig_rx =30;
16819: waveform_sig_rx =242;
16820: waveform_sig_rx =54;
16821: waveform_sig_rx =280;
16822: waveform_sig_rx =127;
16823: waveform_sig_rx =208;
16824: waveform_sig_rx =191;
16825: waveform_sig_rx =77;
16826: waveform_sig_rx =402;
16827: waveform_sig_rx =-8;
16828: waveform_sig_rx =269;
16829: waveform_sig_rx =385;
16830: waveform_sig_rx =-36;
16831: waveform_sig_rx =367;
16832: waveform_sig_rx =382;
16833: waveform_sig_rx =5;
16834: waveform_sig_rx =344;
16835: waveform_sig_rx =417;
16836: waveform_sig_rx =61;
16837: waveform_sig_rx =333;
16838: waveform_sig_rx =422;
16839: waveform_sig_rx =163;
16840: waveform_sig_rx =224;
16841: waveform_sig_rx =491;
16842: waveform_sig_rx =232;
16843: waveform_sig_rx =276;
16844: waveform_sig_rx =323;
16845: waveform_sig_rx =493;
16846: waveform_sig_rx =155;
16847: waveform_sig_rx =314;
16848: waveform_sig_rx =550;
16849: waveform_sig_rx =164;
16850: waveform_sig_rx =306;
16851: waveform_sig_rx =577;
16852: waveform_sig_rx =273;
16853: waveform_sig_rx =291;
16854: waveform_sig_rx =534;
16855: waveform_sig_rx =380;
16856: waveform_sig_rx =314;
16857: waveform_sig_rx =452;
16858: waveform_sig_rx =549;
16859: waveform_sig_rx =310;
16860: waveform_sig_rx =470;
16861: waveform_sig_rx =407;
16862: waveform_sig_rx =512;
16863: waveform_sig_rx =379;
16864: waveform_sig_rx =547;
16865: waveform_sig_rx =384;
16866: waveform_sig_rx =437;
16867: waveform_sig_rx =682;
16868: waveform_sig_rx =199;
16869: waveform_sig_rx =619;
16870: waveform_sig_rx =585;
16871: waveform_sig_rx =264;
16872: waveform_sig_rx =668;
16873: waveform_sig_rx =615;
16874: waveform_sig_rx =270;
16875: waveform_sig_rx =641;
16876: waveform_sig_rx =646;
16877: waveform_sig_rx =319;
16878: waveform_sig_rx =623;
16879: waveform_sig_rx =646;
16880: waveform_sig_rx =463;
16881: waveform_sig_rx =499;
16882: waveform_sig_rx =692;
16883: waveform_sig_rx =562;
16884: waveform_sig_rx =466;
16885: waveform_sig_rx =612;
16886: waveform_sig_rx =768;
16887: waveform_sig_rx =357;
16888: waveform_sig_rx =695;
16889: waveform_sig_rx =766;
16890: waveform_sig_rx =437;
16891: waveform_sig_rx =653;
16892: waveform_sig_rx =763;
16893: waveform_sig_rx =604;
16894: waveform_sig_rx =541;
16895: waveform_sig_rx =763;
16896: waveform_sig_rx =710;
16897: waveform_sig_rx =510;
16898: waveform_sig_rx =731;
16899: waveform_sig_rx =810;
16900: waveform_sig_rx =489;
16901: waveform_sig_rx =768;
16902: waveform_sig_rx =648;
16903: waveform_sig_rx =732;
16904: waveform_sig_rx =679;
16905: waveform_sig_rx =792;
16906: waveform_sig_rx =581;
16907: waveform_sig_rx =735;
16908: waveform_sig_rx =864;
16909: waveform_sig_rx =461;
16910: waveform_sig_rx =904;
16911: waveform_sig_rx =768;
16912: waveform_sig_rx =545;
16913: waveform_sig_rx =923;
16914: waveform_sig_rx =806;
16915: waveform_sig_rx =558;
16916: waveform_sig_rx =871;
16917: waveform_sig_rx =873;
16918: waveform_sig_rx =621;
16919: waveform_sig_rx =829;
16920: waveform_sig_rx =893;
16921: waveform_sig_rx =718;
16922: waveform_sig_rx =665;
16923: waveform_sig_rx =1012;
16924: waveform_sig_rx =784;
16925: waveform_sig_rx =683;
16926: waveform_sig_rx =946;
16927: waveform_sig_rx =928;
16928: waveform_sig_rx =633;
16929: waveform_sig_rx =973;
16930: waveform_sig_rx =898;
16931: waveform_sig_rx =746;
16932: waveform_sig_rx =840;
16933: waveform_sig_rx =950;
16934: waveform_sig_rx =841;
16935: waveform_sig_rx =705;
16936: waveform_sig_rx =1017;
16937: waveform_sig_rx =912;
16938: waveform_sig_rx =698;
16939: waveform_sig_rx =1017;
16940: waveform_sig_rx =999;
16941: waveform_sig_rx =703;
16942: waveform_sig_rx =1029;
16943: waveform_sig_rx =823;
16944: waveform_sig_rx =969;
16945: waveform_sig_rx =905;
16946: waveform_sig_rx =974;
16947: waveform_sig_rx =812;
16948: waveform_sig_rx =1002;
16949: waveform_sig_rx =1009;
16950: waveform_sig_rx =726;
16951: waveform_sig_rx =1119;
16952: waveform_sig_rx =923;
16953: waveform_sig_rx =794;
16954: waveform_sig_rx =1079;
16955: waveform_sig_rx =1006;
16956: waveform_sig_rx =776;
16957: waveform_sig_rx =1045;
16958: waveform_sig_rx =1095;
16959: waveform_sig_rx =786;
16960: waveform_sig_rx =1037;
16961: waveform_sig_rx =1121;
16962: waveform_sig_rx =855;
16963: waveform_sig_rx =900;
16964: waveform_sig_rx =1198;
16965: waveform_sig_rx =905;
16966: waveform_sig_rx =899;
16967: waveform_sig_rx =1107;
16968: waveform_sig_rx =1057;
16969: waveform_sig_rx =852;
16970: waveform_sig_rx =1106;
16971: waveform_sig_rx =1074;
16972: waveform_sig_rx =944;
16973: waveform_sig_rx =975;
16974: waveform_sig_rx =1183;
16975: waveform_sig_rx =1006;
16976: waveform_sig_rx =842;
16977: waveform_sig_rx =1256;
16978: waveform_sig_rx =1002;
16979: waveform_sig_rx =857;
16980: waveform_sig_rx =1227;
16981: waveform_sig_rx =1080;
16982: waveform_sig_rx =922;
16983: waveform_sig_rx =1196;
16984: waveform_sig_rx =927;
16985: waveform_sig_rx =1161;
16986: waveform_sig_rx =1005;
16987: waveform_sig_rx =1120;
16988: waveform_sig_rx =956;
16989: waveform_sig_rx =1103;
16990: waveform_sig_rx =1162;
16991: waveform_sig_rx =872;
16992: waveform_sig_rx =1215;
16993: waveform_sig_rx =1086;
16994: waveform_sig_rx =948;
16995: waveform_sig_rx =1189;
16996: waveform_sig_rx =1170;
16997: waveform_sig_rx =881;
16998: waveform_sig_rx =1192;
16999: waveform_sig_rx =1244;
17000: waveform_sig_rx =850;
17001: waveform_sig_rx =1208;
17002: waveform_sig_rx =1259;
17003: waveform_sig_rx =920;
17004: waveform_sig_rx =1114;
17005: waveform_sig_rx =1272;
17006: waveform_sig_rx =1007;
17007: waveform_sig_rx =1102;
17008: waveform_sig_rx =1161;
17009: waveform_sig_rx =1199;
17010: waveform_sig_rx =957;
17011: waveform_sig_rx =1170;
17012: waveform_sig_rx =1246;
17013: waveform_sig_rx =981;
17014: waveform_sig_rx =1084;
17015: waveform_sig_rx =1330;
17016: waveform_sig_rx =1012;
17017: waveform_sig_rx =998;
17018: waveform_sig_rx =1334;
17019: waveform_sig_rx =1044;
17020: waveform_sig_rx =997;
17021: waveform_sig_rx =1277;
17022: waveform_sig_rx =1141;
17023: waveform_sig_rx =1027;
17024: waveform_sig_rx =1242;
17025: waveform_sig_rx =1012;
17026: waveform_sig_rx =1263;
17027: waveform_sig_rx =1043;
17028: waveform_sig_rx =1230;
17029: waveform_sig_rx =1043;
17030: waveform_sig_rx =1168;
17031: waveform_sig_rx =1258;
17032: waveform_sig_rx =926;
17033: waveform_sig_rx =1290;
17034: waveform_sig_rx =1194;
17035: waveform_sig_rx =950;
17036: waveform_sig_rx =1305;
17037: waveform_sig_rx =1230;
17038: waveform_sig_rx =857;
17039: waveform_sig_rx =1329;
17040: waveform_sig_rx =1230;
17041: waveform_sig_rx =900;
17042: waveform_sig_rx =1319;
17043: waveform_sig_rx =1213;
17044: waveform_sig_rx =998;
17045: waveform_sig_rx =1171;
17046: waveform_sig_rx =1259;
17047: waveform_sig_rx =1107;
17048: waveform_sig_rx =1082;
17049: waveform_sig_rx =1184;
17050: waveform_sig_rx =1267;
17051: waveform_sig_rx =922;
17052: waveform_sig_rx =1260;
17053: waveform_sig_rx =1263;
17054: waveform_sig_rx =985;
17055: waveform_sig_rx =1174;
17056: waveform_sig_rx =1334;
17057: waveform_sig_rx =1023;
17058: waveform_sig_rx =1079;
17059: waveform_sig_rx =1340;
17060: waveform_sig_rx =1054;
17061: waveform_sig_rx =1065;
17062: waveform_sig_rx =1266;
17063: waveform_sig_rx =1171;
17064: waveform_sig_rx =1057;
17065: waveform_sig_rx =1213;
17066: waveform_sig_rx =1062;
17067: waveform_sig_rx =1282;
17068: waveform_sig_rx =1033;
17069: waveform_sig_rx =1267;
17070: waveform_sig_rx =994;
17071: waveform_sig_rx =1174;
17072: waveform_sig_rx =1279;
17073: waveform_sig_rx =875;
17074: waveform_sig_rx =1345;
17075: waveform_sig_rx =1161;
17076: waveform_sig_rx =891;
17077: waveform_sig_rx =1396;
17078: waveform_sig_rx =1128;
17079: waveform_sig_rx =889;
17080: waveform_sig_rx =1351;
17081: waveform_sig_rx =1104;
17082: waveform_sig_rx =968;
17083: waveform_sig_rx =1249;
17084: waveform_sig_rx =1182;
17085: waveform_sig_rx =1014;
17086: waveform_sig_rx =1080;
17087: waveform_sig_rx =1264;
17088: waveform_sig_rx =1063;
17089: waveform_sig_rx =1030;
17090: waveform_sig_rx =1209;
17091: waveform_sig_rx =1181;
17092: waveform_sig_rx =903;
17093: waveform_sig_rx =1241;
17094: waveform_sig_rx =1207;
17095: waveform_sig_rx =901;
17096: waveform_sig_rx =1153;
17097: waveform_sig_rx =1250;
17098: waveform_sig_rx =935;
17099: waveform_sig_rx =1075;
17100: waveform_sig_rx =1212;
17101: waveform_sig_rx =1041;
17102: waveform_sig_rx =989;
17103: waveform_sig_rx =1158;
17104: waveform_sig_rx =1189;
17105: waveform_sig_rx =911;
17106: waveform_sig_rx =1166;
17107: waveform_sig_rx =1025;
17108: waveform_sig_rx =1117;
17109: waveform_sig_rx =1027;
17110: waveform_sig_rx =1172;
17111: waveform_sig_rx =872;
17112: waveform_sig_rx =1202;
17113: waveform_sig_rx =1107;
17114: waveform_sig_rx =809;
17115: waveform_sig_rx =1289;
17116: waveform_sig_rx =974;
17117: waveform_sig_rx =874;
17118: waveform_sig_rx =1270;
17119: waveform_sig_rx =1007;
17120: waveform_sig_rx =853;
17121: waveform_sig_rx =1232;
17122: waveform_sig_rx =1023;
17123: waveform_sig_rx =905;
17124: waveform_sig_rx =1112;
17125: waveform_sig_rx =1074;
17126: waveform_sig_rx =922;
17127: waveform_sig_rx =971;
17128: waveform_sig_rx =1184;
17129: waveform_sig_rx =919;
17130: waveform_sig_rx =909;
17131: waveform_sig_rx =1155;
17132: waveform_sig_rx =1034;
17133: waveform_sig_rx =801;
17134: waveform_sig_rx =1170;
17135: waveform_sig_rx =1025;
17136: waveform_sig_rx =841;
17137: waveform_sig_rx =1057;
17138: waveform_sig_rx =1075;
17139: waveform_sig_rx =880;
17140: waveform_sig_rx =909;
17141: waveform_sig_rx =1089;
17142: waveform_sig_rx =954;
17143: waveform_sig_rx =796;
17144: waveform_sig_rx =1108;
17145: waveform_sig_rx =1021;
17146: waveform_sig_rx =752;
17147: waveform_sig_rx =1121;
17148: waveform_sig_rx =811;
17149: waveform_sig_rx =1004;
17150: waveform_sig_rx =930;
17151: waveform_sig_rx =975;
17152: waveform_sig_rx =776;
17153: waveform_sig_rx =1056;
17154: waveform_sig_rx =920;
17155: waveform_sig_rx =715;
17156: waveform_sig_rx =1120;
17157: waveform_sig_rx =818;
17158: waveform_sig_rx =742;
17159: waveform_sig_rx =1098;
17160: waveform_sig_rx =819;
17161: waveform_sig_rx =727;
17162: waveform_sig_rx =1035;
17163: waveform_sig_rx =837;
17164: waveform_sig_rx =756;
17165: waveform_sig_rx =904;
17166: waveform_sig_rx =964;
17167: waveform_sig_rx =701;
17168: waveform_sig_rx =805;
17169: waveform_sig_rx =1059;
17170: waveform_sig_rx =664;
17171: waveform_sig_rx =799;
17172: waveform_sig_rx =970;
17173: waveform_sig_rx =783;
17174: waveform_sig_rx =702;
17175: waveform_sig_rx =932;
17176: waveform_sig_rx =829;
17177: waveform_sig_rx =684;
17178: waveform_sig_rx =797;
17179: waveform_sig_rx =921;
17180: waveform_sig_rx =667;
17181: waveform_sig_rx =695;
17182: waveform_sig_rx =955;
17183: waveform_sig_rx =693;
17184: waveform_sig_rx =610;
17185: waveform_sig_rx =946;
17186: waveform_sig_rx =743;
17187: waveform_sig_rx =590;
17188: waveform_sig_rx =888;
17189: waveform_sig_rx =575;
17190: waveform_sig_rx =844;
17191: waveform_sig_rx =663;
17192: waveform_sig_rx =760;
17193: waveform_sig_rx =577;
17194: waveform_sig_rx =828;
17195: waveform_sig_rx =688;
17196: waveform_sig_rx =540;
17197: waveform_sig_rx =869;
17198: waveform_sig_rx =611;
17199: waveform_sig_rx =564;
17200: waveform_sig_rx =840;
17201: waveform_sig_rx =644;
17202: waveform_sig_rx =491;
17203: waveform_sig_rx =799;
17204: waveform_sig_rx =670;
17205: waveform_sig_rx =463;
17206: waveform_sig_rx =723;
17207: waveform_sig_rx =758;
17208: waveform_sig_rx =373;
17209: waveform_sig_rx =668;
17210: waveform_sig_rx =732;
17211: waveform_sig_rx =420;
17212: waveform_sig_rx =620;
17213: waveform_sig_rx =641;
17214: waveform_sig_rx =601;
17215: waveform_sig_rx =437;
17216: waveform_sig_rx =669;
17217: waveform_sig_rx =651;
17218: waveform_sig_rx =366;
17219: waveform_sig_rx =605;
17220: waveform_sig_rx =688;
17221: waveform_sig_rx =395;
17222: waveform_sig_rx =481;
17223: waveform_sig_rx =687;
17224: waveform_sig_rx =428;
17225: waveform_sig_rx =385;
17226: waveform_sig_rx =721;
17227: waveform_sig_rx =438;
17228: waveform_sig_rx =400;
17229: waveform_sig_rx =619;
17230: waveform_sig_rx =303;
17231: waveform_sig_rx =639;
17232: waveform_sig_rx =361;
17233: waveform_sig_rx =542;
17234: waveform_sig_rx =337;
17235: waveform_sig_rx =512;
17236: waveform_sig_rx =461;
17237: waveform_sig_rx =271;
17238: waveform_sig_rx =573;
17239: waveform_sig_rx =389;
17240: waveform_sig_rx =217;
17241: waveform_sig_rx =634;
17242: waveform_sig_rx =371;
17243: waveform_sig_rx =159;
17244: waveform_sig_rx =648;
17245: waveform_sig_rx =326;
17246: waveform_sig_rx =210;
17247: waveform_sig_rx =521;
17248: waveform_sig_rx =402;
17249: waveform_sig_rx =174;
17250: waveform_sig_rx =419;
17251: waveform_sig_rx =432;
17252: waveform_sig_rx =229;
17253: waveform_sig_rx =292;
17254: waveform_sig_rx =395;
17255: waveform_sig_rx =354;
17256: waveform_sig_rx =126;
17257: waveform_sig_rx =399;
17258: waveform_sig_rx =345;
17259: waveform_sig_rx =78;
17260: waveform_sig_rx =325;
17261: waveform_sig_rx =422;
17262: waveform_sig_rx =57;
17263: waveform_sig_rx =252;
17264: waveform_sig_rx =412;
17265: waveform_sig_rx =72;
17266: waveform_sig_rx =177;
17267: waveform_sig_rx =363;
17268: waveform_sig_rx =162;
17269: waveform_sig_rx =160;
17270: waveform_sig_rx =237;
17271: waveform_sig_rx =99;
17272: waveform_sig_rx =304;
17273: waveform_sig_rx =50;
17274: waveform_sig_rx =312;
17275: waveform_sig_rx =-25;
17276: waveform_sig_rx =282;
17277: waveform_sig_rx =182;
17278: waveform_sig_rx =-80;
17279: waveform_sig_rx =391;
17280: waveform_sig_rx =51;
17281: waveform_sig_rx =-60;
17282: waveform_sig_rx =402;
17283: waveform_sig_rx =6;
17284: waveform_sig_rx =-68;
17285: waveform_sig_rx =336;
17286: waveform_sig_rx =-27;
17287: waveform_sig_rx =-53;
17288: waveform_sig_rx =210;
17289: waveform_sig_rx =92;
17290: waveform_sig_rx =-111;
17291: waveform_sig_rx =115;
17292: waveform_sig_rx =123;
17293: waveform_sig_rx =-68;
17294: waveform_sig_rx =-50;
17295: waveform_sig_rx =104;
17296: waveform_sig_rx =47;
17297: waveform_sig_rx =-204;
17298: waveform_sig_rx =156;
17299: waveform_sig_rx =20;
17300: waveform_sig_rx =-257;
17301: waveform_sig_rx =94;
17302: waveform_sig_rx =44;
17303: waveform_sig_rx =-230;
17304: waveform_sig_rx =-4;
17305: waveform_sig_rx =5;
17306: waveform_sig_rx =-140;
17307: waveform_sig_rx =-151;
17308: waveform_sig_rx =13;
17309: waveform_sig_rx =-52;
17310: waveform_sig_rx =-234;
17311: waveform_sig_rx =-54;
17312: waveform_sig_rx =-158;
17313: waveform_sig_rx =-89;
17314: waveform_sig_rx =-182;
17315: waveform_sig_rx =-31;
17316: waveform_sig_rx =-383;
17317: waveform_sig_rx =53;
17318: waveform_sig_rx =-210;
17319: waveform_sig_rx =-337;
17320: waveform_sig_rx =82;
17321: waveform_sig_rx =-321;
17322: waveform_sig_rx =-301;
17323: waveform_sig_rx =50;
17324: waveform_sig_rx =-329;
17325: waveform_sig_rx =-364;
17326: waveform_sig_rx =8;
17327: waveform_sig_rx =-343;
17328: waveform_sig_rx =-329;
17329: waveform_sig_rx =-116;
17330: waveform_sig_rx =-242;
17331: waveform_sig_rx =-388;
17332: waveform_sig_rx =-231;
17333: waveform_sig_rx =-143;
17334: waveform_sig_rx =-357;
17335: waveform_sig_rx =-386;
17336: waveform_sig_rx =-103;
17337: waveform_sig_rx =-345;
17338: waveform_sig_rx =-497;
17339: waveform_sig_rx =-81;
17340: waveform_sig_rx =-398;
17341: waveform_sig_rx =-441;
17342: waveform_sig_rx =-220;
17343: waveform_sig_rx =-286;
17344: waveform_sig_rx =-453;
17345: waveform_sig_rx =-380;
17346: waveform_sig_rx =-225;
17347: waveform_sig_rx =-435;
17348: waveform_sig_rx =-494;
17349: waveform_sig_rx =-192;
17350: waveform_sig_rx =-440;
17351: waveform_sig_rx =-510;
17352: waveform_sig_rx =-306;
17353: waveform_sig_rx =-505;
17354: waveform_sig_rx =-360;
17355: waveform_sig_rx =-451;
17356: waveform_sig_rx =-380;
17357: waveform_sig_rx =-624;
17358: waveform_sig_rx =-229;
17359: waveform_sig_rx =-572;
17360: waveform_sig_rx =-568;
17361: waveform_sig_rx =-233;
17362: waveform_sig_rx =-651;
17363: waveform_sig_rx =-530;
17364: waveform_sig_rx =-290;
17365: waveform_sig_rx =-622;
17366: waveform_sig_rx =-600;
17367: waveform_sig_rx =-330;
17368: waveform_sig_rx =-593;
17369: waveform_sig_rx =-624;
17370: waveform_sig_rx =-416;
17371: waveform_sig_rx =-448;
17372: waveform_sig_rx =-734;
17373: waveform_sig_rx =-493;
17374: waveform_sig_rx =-410;
17375: waveform_sig_rx =-715;
17376: waveform_sig_rx =-623;
17377: waveform_sig_rx =-385;
17378: waveform_sig_rx =-701;
17379: waveform_sig_rx =-706;
17380: waveform_sig_rx =-431;
17381: waveform_sig_rx =-673;
17382: waveform_sig_rx =-690;
17383: waveform_sig_rx =-587;
17384: waveform_sig_rx =-519;
17385: waveform_sig_rx =-766;
17386: waveform_sig_rx =-693;
17387: waveform_sig_rx =-455;
17388: waveform_sig_rx =-807;
17389: waveform_sig_rx =-750;
17390: waveform_sig_rx =-449;
17391: waveform_sig_rx =-775;
17392: waveform_sig_rx =-743;
17393: waveform_sig_rx =-608;
17394: waveform_sig_rx =-797;
17395: waveform_sig_rx =-593;
17396: waveform_sig_rx =-736;
17397: waveform_sig_rx =-643;
17398: waveform_sig_rx =-843;
17399: waveform_sig_rx =-522;
17400: waveform_sig_rx =-846;
17401: waveform_sig_rx =-793;
17402: waveform_sig_rx =-569;
17403: waveform_sig_rx =-887;
17404: waveform_sig_rx =-798;
17405: waveform_sig_rx =-598;
17406: waveform_sig_rx =-823;
17407: waveform_sig_rx =-901;
17408: waveform_sig_rx =-559;
17409: waveform_sig_rx =-824;
17410: waveform_sig_rx =-938;
17411: waveform_sig_rx =-633;
17412: waveform_sig_rx =-757;
17413: waveform_sig_rx =-1018;
17414: waveform_sig_rx =-703;
17415: waveform_sig_rx =-735;
17416: waveform_sig_rx =-966;
17417: waveform_sig_rx =-839;
17418: waveform_sig_rx =-696;
17419: waveform_sig_rx =-907;
17420: waveform_sig_rx =-929;
17421: waveform_sig_rx =-718;
17422: waveform_sig_rx =-853;
17423: waveform_sig_rx =-968;
17424: waveform_sig_rx =-821;
17425: waveform_sig_rx =-689;
17426: waveform_sig_rx =-1078;
17427: waveform_sig_rx =-872;
17428: waveform_sig_rx =-671;
17429: waveform_sig_rx =-1076;
17430: waveform_sig_rx =-886;
17431: waveform_sig_rx =-707;
17432: waveform_sig_rx =-1011;
17433: waveform_sig_rx =-898;
17434: waveform_sig_rx =-879;
17435: waveform_sig_rx =-977;
17436: waveform_sig_rx =-814;
17437: waveform_sig_rx =-982;
17438: waveform_sig_rx =-841;
17439: waveform_sig_rx =-1067;
17440: waveform_sig_rx =-759;
17441: waveform_sig_rx =-1033;
17442: waveform_sig_rx =-1012;
17443: waveform_sig_rx =-773;
17444: waveform_sig_rx =-1059;
17445: waveform_sig_rx =-1038;
17446: waveform_sig_rx =-760;
17447: waveform_sig_rx =-1045;
17448: waveform_sig_rx =-1152;
17449: waveform_sig_rx =-723;
17450: waveform_sig_rx =-1074;
17451: waveform_sig_rx =-1126;
17452: waveform_sig_rx =-792;
17453: waveform_sig_rx =-1011;
17454: waveform_sig_rx =-1159;
17455: waveform_sig_rx =-854;
17456: waveform_sig_rx =-968;
17457: waveform_sig_rx =-1102;
17458: waveform_sig_rx =-1039;
17459: waveform_sig_rx =-887;
17460: waveform_sig_rx =-1051;
17461: waveform_sig_rx =-1153;
17462: waveform_sig_rx =-865;
17463: waveform_sig_rx =-1029;
17464: waveform_sig_rx =-1207;
17465: waveform_sig_rx =-921;
17466: waveform_sig_rx =-929;
17467: waveform_sig_rx =-1265;
17468: waveform_sig_rx =-959;
17469: waveform_sig_rx =-940;
17470: waveform_sig_rx =-1225;
17471: waveform_sig_rx =-1070;
17472: waveform_sig_rx =-922;
17473: waveform_sig_rx =-1136;
17474: waveform_sig_rx =-1090;
17475: waveform_sig_rx =-1059;
17476: waveform_sig_rx =-1126;
17477: waveform_sig_rx =-1022;
17478: waveform_sig_rx =-1135;
17479: waveform_sig_rx =-995;
17480: waveform_sig_rx =-1260;
17481: waveform_sig_rx =-914;
17482: waveform_sig_rx =-1198;
17483: waveform_sig_rx =-1175;
17484: waveform_sig_rx =-911;
17485: waveform_sig_rx =-1211;
17486: waveform_sig_rx =-1192;
17487: waveform_sig_rx =-848;
17488: waveform_sig_rx =-1242;
17489: waveform_sig_rx =-1268;
17490: waveform_sig_rx =-794;
17491: waveform_sig_rx =-1312;
17492: waveform_sig_rx =-1162;
17493: waveform_sig_rx =-941;
17494: waveform_sig_rx =-1214;
17495: waveform_sig_rx =-1232;
17496: waveform_sig_rx =-1061;
17497: waveform_sig_rx =-1082;
17498: waveform_sig_rx =-1206;
17499: waveform_sig_rx =-1228;
17500: waveform_sig_rx =-947;
17501: waveform_sig_rx =-1239;
17502: waveform_sig_rx =-1272;
17503: waveform_sig_rx =-921;
17504: waveform_sig_rx =-1211;
17505: waveform_sig_rx =-1259;
17506: waveform_sig_rx =-1010;
17507: waveform_sig_rx =-1079;
17508: waveform_sig_rx =-1323;
17509: waveform_sig_rx =-1065;
17510: waveform_sig_rx =-1042;
17511: waveform_sig_rx =-1288;
17512: waveform_sig_rx =-1151;
17513: waveform_sig_rx =-1024;
17514: waveform_sig_rx =-1239;
17515: waveform_sig_rx =-1158;
17516: waveform_sig_rx =-1155;
17517: waveform_sig_rx =-1152;
17518: waveform_sig_rx =-1114;
17519: waveform_sig_rx =-1179;
17520: waveform_sig_rx =-1082;
17521: waveform_sig_rx =-1358;
17522: waveform_sig_rx =-923;
17523: waveform_sig_rx =-1295;
17524: waveform_sig_rx =-1251;
17525: waveform_sig_rx =-917;
17526: waveform_sig_rx =-1381;
17527: waveform_sig_rx =-1196;
17528: waveform_sig_rx =-919;
17529: waveform_sig_rx =-1395;
17530: waveform_sig_rx =-1176;
17531: waveform_sig_rx =-959;
17532: waveform_sig_rx =-1319;
17533: waveform_sig_rx =-1160;
17534: waveform_sig_rx =-1073;
17535: waveform_sig_rx =-1157;
17536: waveform_sig_rx =-1326;
17537: waveform_sig_rx =-1085;
17538: waveform_sig_rx =-1075;
17539: waveform_sig_rx =-1306;
17540: waveform_sig_rx =-1189;
17541: waveform_sig_rx =-978;
17542: waveform_sig_rx =-1292;
17543: waveform_sig_rx =-1237;
17544: waveform_sig_rx =-979;
17545: waveform_sig_rx =-1231;
17546: waveform_sig_rx =-1265;
17547: waveform_sig_rx =-1024;
17548: waveform_sig_rx =-1113;
17549: waveform_sig_rx =-1313;
17550: waveform_sig_rx =-1089;
17551: waveform_sig_rx =-1068;
17552: waveform_sig_rx =-1256;
17553: waveform_sig_rx =-1208;
17554: waveform_sig_rx =-985;
17555: waveform_sig_rx =-1221;
17556: waveform_sig_rx =-1184;
17557: waveform_sig_rx =-1085;
17558: waveform_sig_rx =-1182;
17559: waveform_sig_rx =-1143;
17560: waveform_sig_rx =-1130;
17561: waveform_sig_rx =-1147;
17562: waveform_sig_rx =-1297;
17563: waveform_sig_rx =-890;
17564: waveform_sig_rx =-1365;
17565: waveform_sig_rx =-1121;
17566: waveform_sig_rx =-945;
17567: waveform_sig_rx =-1367;
17568: waveform_sig_rx =-1077;
17569: waveform_sig_rx =-992;
17570: waveform_sig_rx =-1281;
17571: waveform_sig_rx =-1150;
17572: waveform_sig_rx =-962;
17573: waveform_sig_rx =-1240;
17574: waveform_sig_rx =-1193;
17575: waveform_sig_rx =-984;
17576: waveform_sig_rx =-1096;
17577: waveform_sig_rx =-1315;
17578: waveform_sig_rx =-970;
17579: waveform_sig_rx =-1073;
17580: waveform_sig_rx =-1236;
17581: waveform_sig_rx =-1125;
17582: waveform_sig_rx =-949;
17583: waveform_sig_rx =-1231;
17584: waveform_sig_rx =-1165;
17585: waveform_sig_rx =-897;
17586: waveform_sig_rx =-1206;
17587: waveform_sig_rx =-1157;
17588: waveform_sig_rx =-975;
17589: waveform_sig_rx =-1064;
17590: waveform_sig_rx =-1181;
17591: waveform_sig_rx =-1061;
17592: waveform_sig_rx =-933;
17593: waveform_sig_rx =-1213;
17594: waveform_sig_rx =-1148;
17595: waveform_sig_rx =-804;
17596: waveform_sig_rx =-1261;
17597: waveform_sig_rx =-1041;
17598: waveform_sig_rx =-1018;
17599: waveform_sig_rx =-1153;
17600: waveform_sig_rx =-951;
17601: waveform_sig_rx =-1080;
17602: waveform_sig_rx =-1063;
17603: waveform_sig_rx =-1131;
17604: waveform_sig_rx =-851;
17605: waveform_sig_rx =-1229;
17606: waveform_sig_rx =-1012;
17607: waveform_sig_rx =-909;
17608: waveform_sig_rx =-1205;
17609: waveform_sig_rx =-1000;
17610: waveform_sig_rx =-842;
17611: waveform_sig_rx =-1193;
17612: waveform_sig_rx =-1060;
17613: waveform_sig_rx =-834;
17614: waveform_sig_rx =-1148;
17615: waveform_sig_rx =-1057;
17616: waveform_sig_rx =-878;
17617: waveform_sig_rx =-974;
17618: waveform_sig_rx =-1212;
17619: waveform_sig_rx =-809;
17620: waveform_sig_rx =-956;
17621: waveform_sig_rx =-1140;
17622: waveform_sig_rx =-921;
17623: waveform_sig_rx =-854;
17624: waveform_sig_rx =-1087;
17625: waveform_sig_rx =-968;
17626: waveform_sig_rx =-850;
17627: waveform_sig_rx =-1010;
17628: waveform_sig_rx =-1052;
17629: waveform_sig_rx =-849;
17630: waveform_sig_rx =-855;
17631: waveform_sig_rx =-1134;
17632: waveform_sig_rx =-848;
17633: waveform_sig_rx =-783;
17634: waveform_sig_rx =-1132;
17635: waveform_sig_rx =-886;
17636: waveform_sig_rx =-717;
17637: waveform_sig_rx =-1108;
17638: waveform_sig_rx =-822;
17639: waveform_sig_rx =-954;
17640: waveform_sig_rx =-953;
17641: waveform_sig_rx =-815;
17642: waveform_sig_rx =-987;
17643: waveform_sig_rx =-846;
17644: waveform_sig_rx =-1003;
17645: waveform_sig_rx =-704;
17646: waveform_sig_rx =-1031;
17647: waveform_sig_rx =-889;
17648: waveform_sig_rx =-713;
17649: waveform_sig_rx =-1042;
17650: waveform_sig_rx =-847;
17651: waveform_sig_rx =-665;
17652: waveform_sig_rx =-1035;
17653: waveform_sig_rx =-877;
17654: waveform_sig_rx =-637;
17655: waveform_sig_rx =-987;
17656: waveform_sig_rx =-873;
17657: waveform_sig_rx =-638;
17658: waveform_sig_rx =-845;
17659: waveform_sig_rx =-991;
17660: waveform_sig_rx =-561;
17661: waveform_sig_rx =-840;
17662: waveform_sig_rx =-869;
17663: waveform_sig_rx =-731;
17664: waveform_sig_rx =-702;
17665: waveform_sig_rx =-814;
17666: waveform_sig_rx =-839;
17667: waveform_sig_rx =-608;
17668: waveform_sig_rx =-779;
17669: waveform_sig_rx =-906;
17670: waveform_sig_rx =-565;
17671: waveform_sig_rx =-714;
17672: waveform_sig_rx =-915;
17673: waveform_sig_rx =-578;
17674: waveform_sig_rx =-654;
17675: waveform_sig_rx =-872;
17676: waveform_sig_rx =-663;
17677: waveform_sig_rx =-570;
17678: waveform_sig_rx =-854;
17679: waveform_sig_rx =-604;
17680: waveform_sig_rx =-753;
17681: waveform_sig_rx =-660;
17682: waveform_sig_rx =-615;
17683: waveform_sig_rx =-719;
17684: waveform_sig_rx =-603;
17685: waveform_sig_rx =-800;
17686: waveform_sig_rx =-455;
17687: waveform_sig_rx =-799;
17688: waveform_sig_rx =-668;
17689: waveform_sig_rx =-454;
17690: waveform_sig_rx =-825;
17691: waveform_sig_rx =-629;
17692: waveform_sig_rx =-401;
17693: waveform_sig_rx =-841;
17694: waveform_sig_rx =-618;
17695: waveform_sig_rx =-377;
17696: waveform_sig_rx =-824;
17697: waveform_sig_rx =-588;
17698: waveform_sig_rx =-438;
17699: waveform_sig_rx =-656;
17700: waveform_sig_rx =-696;
17701: waveform_sig_rx =-406;
17702: waveform_sig_rx =-603;
17703: waveform_sig_rx =-598;
17704: waveform_sig_rx =-565;
17705: waveform_sig_rx =-392;
17706: waveform_sig_rx =-631;
17707: waveform_sig_rx =-603;
17708: waveform_sig_rx =-304;
17709: waveform_sig_rx =-611;
17710: waveform_sig_rx =-631;
17711: waveform_sig_rx =-301;
17712: waveform_sig_rx =-514;
17713: waveform_sig_rx =-626;
17714: waveform_sig_rx =-338;
17715: waveform_sig_rx =-415;
17716: waveform_sig_rx =-607;
17717: waveform_sig_rx =-413;
17718: waveform_sig_rx =-308;
17719: waveform_sig_rx =-592;
17720: waveform_sig_rx =-370;
17721: waveform_sig_rx =-493;
17722: waveform_sig_rx =-362;
17723: waveform_sig_rx =-422;
17724: waveform_sig_rx =-407;
17725: waveform_sig_rx =-364;
17726: waveform_sig_rx =-560;
17727: waveform_sig_rx =-135;
17728: waveform_sig_rx =-592;
17729: waveform_sig_rx =-352;
17730: waveform_sig_rx =-162;
17731: waveform_sig_rx =-616;
17732: waveform_sig_rx =-256;
17733: waveform_sig_rx =-154;
17734: waveform_sig_rx =-590;
17735: waveform_sig_rx =-274;
17736: waveform_sig_rx =-143;
17737: waveform_sig_rx =-505;
17738: waveform_sig_rx =-291;
17739: waveform_sig_rx =-192;
17740: waveform_sig_rx =-352;
17741: waveform_sig_rx =-410;
17742: waveform_sig_rx =-135;
17743: waveform_sig_rx =-291;
17744: waveform_sig_rx =-328;
17745: waveform_sig_rx =-268;
17746: waveform_sig_rx =-77;
17747: waveform_sig_rx =-400;
17748: waveform_sig_rx =-295;
17749: waveform_sig_rx =-14;
17750: waveform_sig_rx =-389;
17751: waveform_sig_rx =-276;
17752: waveform_sig_rx =-41;
17753: waveform_sig_rx =-272;
17754: waveform_sig_rx =-306;
17755: waveform_sig_rx =-102;
17756: waveform_sig_rx =-132;
17757: waveform_sig_rx =-293;
17758: waveform_sig_rx =-156;
17759: waveform_sig_rx =12;
17760: waveform_sig_rx =-305;
17761: waveform_sig_rx =-99;
17762: waveform_sig_rx =-160;
17763: waveform_sig_rx =-125;
17764: waveform_sig_rx =-144;
17765: waveform_sig_rx =-68;
17766: waveform_sig_rx =-142;
17767: waveform_sig_rx =-200;
17768: waveform_sig_rx =143;
17769: waveform_sig_rx =-352;
17770: waveform_sig_rx =-5;
17771: waveform_sig_rx =70;
17772: waveform_sig_rx =-326;
17773: waveform_sig_rx =64;
17774: waveform_sig_rx =83;
17775: waveform_sig_rx =-276;
17776: waveform_sig_rx =30;
17777: waveform_sig_rx =97;
17778: waveform_sig_rx =-196;
17779: waveform_sig_rx =-4;
17780: waveform_sig_rx =84;
17781: waveform_sig_rx =-48;
17782: waveform_sig_rx =-139;
17783: waveform_sig_rx =165;
17784: waveform_sig_rx =25;
17785: waveform_sig_rx =-112;
17786: waveform_sig_rx =52;
17787: waveform_sig_rx =214;
17788: waveform_sig_rx =-157;
17789: waveform_sig_rx =97;
17790: waveform_sig_rx =235;
17791: waveform_sig_rx =-54;
17792: waveform_sig_rx =64;
17793: waveform_sig_rx =217;
17794: waveform_sig_rx =102;
17795: waveform_sig_rx =-33;
17796: waveform_sig_rx =198;
17797: waveform_sig_rx =205;
17798: waveform_sig_rx =-46;
17799: waveform_sig_rx =152;
17800: waveform_sig_rx =300;
17801: waveform_sig_rx =-49;
17802: waveform_sig_rx =233;
17803: waveform_sig_rx =127;
17804: waveform_sig_rx =163;
17805: waveform_sig_rx =157;
17806: waveform_sig_rx =210;
17807: waveform_sig_rx =120;
17808: waveform_sig_rx =146;
17809: waveform_sig_rx =382;
17810: waveform_sig_rx =-48;
17811: waveform_sig_rx =341;
17812: waveform_sig_rx =304;
17813: waveform_sig_rx =14;
17814: waveform_sig_rx =363;
17815: waveform_sig_rx =347;
17816: waveform_sig_rx =57;
17817: waveform_sig_rx =309;
17818: waveform_sig_rx =415;
17819: waveform_sig_rx =120;
17820: waveform_sig_rx =282;
17821: waveform_sig_rx =408;
17822: waveform_sig_rx =236;
17823: waveform_sig_rx =132;
17824: waveform_sig_rx =506;
17825: waveform_sig_rx =283;
17826: waveform_sig_rx =168;
17827: waveform_sig_rx =413;
17828: waveform_sig_rx =428;
17829: waveform_sig_rx =175;
17830: waveform_sig_rx =410;
17831: waveform_sig_rx =446;
17832: waveform_sig_rx =283;
17833: waveform_sig_rx =306;
17834: waveform_sig_rx =488;
17835: waveform_sig_rx =393;
17836: waveform_sig_rx =213;
17837: waveform_sig_rx =544;
17838: waveform_sig_rx =460;
17839: waveform_sig_rx =219;
17840: waveform_sig_rx =489;
17841: waveform_sig_rx =548;
17842: waveform_sig_rx =242;
17843: waveform_sig_rx =548;
17844: waveform_sig_rx =388;
17845: waveform_sig_rx =460;
17846: waveform_sig_rx =468;
17847: waveform_sig_rx =481;
17848: waveform_sig_rx =406;
17849: waveform_sig_rx =456;
17850: waveform_sig_rx =617;
17851: waveform_sig_rx =285;
17852: waveform_sig_rx =598;
17853: waveform_sig_rx =541;
17854: waveform_sig_rx =351;
17855: waveform_sig_rx =567;
17856: waveform_sig_rx =657;
17857: waveform_sig_rx =332;
17858: waveform_sig_rx =557;
17859: waveform_sig_rx =730;
17860: waveform_sig_rx =307;
17861: waveform_sig_rx =587;
17862: waveform_sig_rx =696;
17863: waveform_sig_rx =438;
17864: waveform_sig_rx =441;
17865: waveform_sig_rx =754;
17866: waveform_sig_rx =520;
17867: waveform_sig_rx =493;
17868: waveform_sig_rx =656;
17869: waveform_sig_rx =695;
17870: waveform_sig_rx =429;
17871: waveform_sig_rx =644;
17872: waveform_sig_rx =725;
17873: waveform_sig_rx =544;
17874: waveform_sig_rx =555;
17875: waveform_sig_rx =810;
17876: waveform_sig_rx =654;
17877: waveform_sig_rx =440;
17878: waveform_sig_rx =853;
17879: waveform_sig_rx =660;
17880: waveform_sig_rx =491;
17881: waveform_sig_rx =807;
17882: waveform_sig_rx =737;
17883: waveform_sig_rx =546;
17884: waveform_sig_rx =772;
17885: waveform_sig_rx =595;
17886: waveform_sig_rx =786;
17887: waveform_sig_rx =672;
17888: waveform_sig_rx =745;
17889: waveform_sig_rx =677;
17890: waveform_sig_rx =661;
17891: waveform_sig_rx =883;
17892: waveform_sig_rx =531;
17893: waveform_sig_rx =806;
17894: waveform_sig_rx =829;
17895: waveform_sig_rx =551;
17896: waveform_sig_rx =832;
17897: waveform_sig_rx =907;
17898: waveform_sig_rx =515;
17899: waveform_sig_rx =832;
17900: waveform_sig_rx =947;
17901: waveform_sig_rx =531;
17902: waveform_sig_rx =849;
17903: waveform_sig_rx =926;
17904: waveform_sig_rx =658;
17905: waveform_sig_rx =725;
17906: waveform_sig_rx =972;
17907: waveform_sig_rx =744;
17908: waveform_sig_rx =753;
17909: waveform_sig_rx =840;
17910: waveform_sig_rx =943;
17911: waveform_sig_rx =674;
17912: waveform_sig_rx =850;
17913: waveform_sig_rx =981;
17914: waveform_sig_rx =709;
17915: waveform_sig_rx =777;
17916: waveform_sig_rx =1058;
17917: waveform_sig_rx =788;
17918: waveform_sig_rx =712;
17919: waveform_sig_rx =1069;
17920: waveform_sig_rx =833;
17921: waveform_sig_rx =751;
17922: waveform_sig_rx =969;
17923: waveform_sig_rx =939;
17924: waveform_sig_rx =775;
17925: waveform_sig_rx =945;
17926: waveform_sig_rx =826;
17927: waveform_sig_rx =978;
17928: waveform_sig_rx =837;
17929: waveform_sig_rx =987;
17930: waveform_sig_rx =854;
17931: waveform_sig_rx =884;
17932: waveform_sig_rx =1103;
17933: waveform_sig_rx =694;
17934: waveform_sig_rx =1036;
17935: waveform_sig_rx =1037;
17936: waveform_sig_rx =718;
17937: waveform_sig_rx =1080;
17938: waveform_sig_rx =1093;
17939: waveform_sig_rx =688;
17940: waveform_sig_rx =1095;
17941: waveform_sig_rx =1118;
17942: waveform_sig_rx =732;
17943: waveform_sig_rx =1108;
17944: waveform_sig_rx =1052;
17945: waveform_sig_rx =878;
17946: waveform_sig_rx =948;
17947: waveform_sig_rx =1099;
17948: waveform_sig_rx =980;
17949: waveform_sig_rx =897;
17950: waveform_sig_rx =1035;
17951: waveform_sig_rx =1158;
17952: waveform_sig_rx =784;
17953: waveform_sig_rx =1099;
17954: waveform_sig_rx =1161;
17955: waveform_sig_rx =850;
17956: waveform_sig_rx =1006;
17957: waveform_sig_rx =1175;
17958: waveform_sig_rx =935;
17959: waveform_sig_rx =913;
17960: waveform_sig_rx =1204;
17961: waveform_sig_rx =1019;
17962: waveform_sig_rx =918;
17963: waveform_sig_rx =1121;
17964: waveform_sig_rx =1142;
17965: waveform_sig_rx =911;
17966: waveform_sig_rx =1114;
17967: waveform_sig_rx =999;
17968: waveform_sig_rx =1123;
17969: waveform_sig_rx =987;
17970: waveform_sig_rx =1154;
17971: waveform_sig_rx =964;
17972: waveform_sig_rx =1066;
17973: waveform_sig_rx =1238;
17974: waveform_sig_rx =818;
17975: waveform_sig_rx =1216;
17976: waveform_sig_rx =1154;
17977: waveform_sig_rx =821;
17978: waveform_sig_rx =1288;
17979: waveform_sig_rx =1150;
17980: waveform_sig_rx =831;
17981: waveform_sig_rx =1284;
17982: waveform_sig_rx =1140;
17983: waveform_sig_rx =926;
17984: waveform_sig_rx =1200;
17985: waveform_sig_rx =1154;
17986: waveform_sig_rx =1062;
17987: waveform_sig_rx =974;
17988: waveform_sig_rx =1278;
17989: waveform_sig_rx =1076;
17990: waveform_sig_rx =968;
17991: waveform_sig_rx =1231;
17992: waveform_sig_rx =1184;
17993: waveform_sig_rx =924;
17994: waveform_sig_rx =1228;
17995: waveform_sig_rx =1192;
17996: waveform_sig_rx =989;
17997: waveform_sig_rx =1101;
17998: waveform_sig_rx =1265;
17999: waveform_sig_rx =1033;
18000: waveform_sig_rx =1027;
18001: waveform_sig_rx =1289;
18002: waveform_sig_rx =1106;
18003: waveform_sig_rx =1015;
18004: waveform_sig_rx =1208;
18005: waveform_sig_rx =1237;
18006: waveform_sig_rx =965;
18007: waveform_sig_rx =1183;
18008: waveform_sig_rx =1110;
18009: waveform_sig_rx =1158;
18010: waveform_sig_rx =1092;
18011: waveform_sig_rx =1254;
18012: waveform_sig_rx =963;
18013: waveform_sig_rx =1210;
18014: waveform_sig_rx =1243;
18015: waveform_sig_rx =881;
18016: waveform_sig_rx =1365;
18017: waveform_sig_rx =1115;
18018: waveform_sig_rx =969;
18019: waveform_sig_rx =1314;
18020: waveform_sig_rx =1157;
18021: waveform_sig_rx =958;
18022: waveform_sig_rx =1262;
18023: waveform_sig_rx =1227;
18024: waveform_sig_rx =988;
18025: waveform_sig_rx =1209;
18026: waveform_sig_rx =1258;
18027: waveform_sig_rx =1032;
18028: waveform_sig_rx =1069;
18029: waveform_sig_rx =1351;
18030: waveform_sig_rx =1062;
18031: waveform_sig_rx =1051;
18032: waveform_sig_rx =1243;
18033: waveform_sig_rx =1211;
18034: waveform_sig_rx =958;
18035: waveform_sig_rx =1258;
18036: waveform_sig_rx =1227;
18037: waveform_sig_rx =1000;
18038: waveform_sig_rx =1155;
18039: waveform_sig_rx =1281;
18040: waveform_sig_rx =1085;
18041: waveform_sig_rx =1049;
18042: waveform_sig_rx =1278;
18043: waveform_sig_rx =1171;
18044: waveform_sig_rx =968;
18045: waveform_sig_rx =1268;
18046: waveform_sig_rx =1261;
18047: waveform_sig_rx =946;
18048: waveform_sig_rx =1311;
18049: waveform_sig_rx =1038;
18050: waveform_sig_rx =1202;
18051: waveform_sig_rx =1148;
18052: waveform_sig_rx =1179;
18053: waveform_sig_rx =1035;
18054: waveform_sig_rx =1228;
18055: waveform_sig_rx =1187;
18056: waveform_sig_rx =942;
18057: waveform_sig_rx =1303;
18058: waveform_sig_rx =1116;
18059: waveform_sig_rx =995;
18060: waveform_sig_rx =1289;
18061: waveform_sig_rx =1195;
18062: waveform_sig_rx =919;
18063: waveform_sig_rx =1286;
18064: waveform_sig_rx =1206;
18065: waveform_sig_rx =955;
18066: waveform_sig_rx =1218;
18067: waveform_sig_rx =1235;
18068: waveform_sig_rx =986;
18069: waveform_sig_rx =1060;
18070: waveform_sig_rx =1314;
18071: waveform_sig_rx =1010;
18072: waveform_sig_rx =1034;
18073: waveform_sig_rx =1217;
18074: waveform_sig_rx =1131;
18075: waveform_sig_rx =947;
18076: waveform_sig_rx =1224;
18077: waveform_sig_rx =1150;
18078: waveform_sig_rx =999;
18079: waveform_sig_rx =1074;
18080: waveform_sig_rx =1236;
18081: waveform_sig_rx =1037;
18082: waveform_sig_rx =934;
18083: waveform_sig_rx =1313;
18084: waveform_sig_rx =1054;
18085: waveform_sig_rx =909;
18086: waveform_sig_rx =1278;
18087: waveform_sig_rx =1080;
18088: waveform_sig_rx =960;
18089: waveform_sig_rx =1225;
18090: waveform_sig_rx =920;
18091: waveform_sig_rx =1240;
18092: waveform_sig_rx =990;
18093: waveform_sig_rx =1148;
18094: waveform_sig_rx =990;
18095: waveform_sig_rx =1097;
18096: waveform_sig_rx =1167;
18097: waveform_sig_rx =842;
18098: waveform_sig_rx =1222;
18099: waveform_sig_rx =1065;
18100: waveform_sig_rx =854;
18101: waveform_sig_rx =1253;
18102: waveform_sig_rx =1050;
18103: waveform_sig_rx =851;
18104: waveform_sig_rx =1193;
18105: waveform_sig_rx =1091;
18106: waveform_sig_rx =852;
18107: waveform_sig_rx =1088;
18108: waveform_sig_rx =1157;
18109: waveform_sig_rx =825;
18110: waveform_sig_rx =1013;
18111: waveform_sig_rx =1176;
18112: waveform_sig_rx =861;
18113: waveform_sig_rx =1015;
18114: waveform_sig_rx =1068;
18115: waveform_sig_rx =1065;
18116: waveform_sig_rx =858;
18117: waveform_sig_rx =1051;
18118: waveform_sig_rx =1130;
18119: waveform_sig_rx =812;
18120: waveform_sig_rx =982;
18121: waveform_sig_rx =1172;
18122: waveform_sig_rx =832;
18123: waveform_sig_rx =915;
18124: waveform_sig_rx =1159;
18125: waveform_sig_rx =886;
18126: waveform_sig_rx =853;
18127: waveform_sig_rx =1099;
18128: waveform_sig_rx =968;
18129: waveform_sig_rx =845;
18130: waveform_sig_rx =1043;
18131: waveform_sig_rx =813;
18132: waveform_sig_rx =1068;
18133: waveform_sig_rx =821;
18134: waveform_sig_rx =1045;
18135: waveform_sig_rx =801;
18136: waveform_sig_rx =967;
18137: waveform_sig_rx =1017;
18138: waveform_sig_rx =687;
18139: waveform_sig_rx =1099;
18140: waveform_sig_rx =911;
18141: waveform_sig_rx =691;
18142: waveform_sig_rx =1112;
18143: waveform_sig_rx =903;
18144: waveform_sig_rx =660;
18145: waveform_sig_rx =1073;
18146: waveform_sig_rx =899;
18147: waveform_sig_rx =687;
18148: waveform_sig_rx =991;
18149: waveform_sig_rx =944;
18150: waveform_sig_rx =680;
18151: waveform_sig_rx =865;
18152: waveform_sig_rx =946;
18153: waveform_sig_rx =749;
18154: waveform_sig_rx =799;
18155: waveform_sig_rx =886;
18156: waveform_sig_rx =936;
18157: waveform_sig_rx =606;
18158: waveform_sig_rx =933;
18159: waveform_sig_rx =908;
18160: waveform_sig_rx =572;
18161: waveform_sig_rx =880;
18162: waveform_sig_rx =927;
18163: waveform_sig_rx =645;
18164: waveform_sig_rx =761;
18165: waveform_sig_rx =910;
18166: waveform_sig_rx =733;
18167: waveform_sig_rx =658;
18168: waveform_sig_rx =895;
18169: waveform_sig_rx =789;
18170: waveform_sig_rx =624;
18171: waveform_sig_rx =829;
18172: waveform_sig_rx =645;
18173: waveform_sig_rx =845;
18174: waveform_sig_rx =637;
18175: waveform_sig_rx =854;
18176: waveform_sig_rx =549;
18177: waveform_sig_rx =822;
18178: waveform_sig_rx =795;
18179: waveform_sig_rx =460;
18180: waveform_sig_rx =929;
18181: waveform_sig_rx =666;
18182: waveform_sig_rx =486;
18183: waveform_sig_rx =943;
18184: waveform_sig_rx =617;
18185: waveform_sig_rx =477;
18186: waveform_sig_rx =890;
18187: waveform_sig_rx =606;
18188: waveform_sig_rx =537;
18189: waveform_sig_rx =753;
18190: waveform_sig_rx =682;
18191: waveform_sig_rx =506;
18192: waveform_sig_rx =588;
18193: waveform_sig_rx =748;
18194: waveform_sig_rx =514;
18195: waveform_sig_rx =512;
18196: waveform_sig_rx =707;
18197: waveform_sig_rx =627;
18198: waveform_sig_rx =360;
18199: waveform_sig_rx =745;
18200: waveform_sig_rx =605;
18201: waveform_sig_rx =384;
18202: waveform_sig_rx =636;
18203: waveform_sig_rx =640;
18204: waveform_sig_rx =442;
18205: waveform_sig_rx =500;
18206: waveform_sig_rx =658;
18207: waveform_sig_rx =504;
18208: waveform_sig_rx =387;
18209: waveform_sig_rx =658;
18210: waveform_sig_rx =531;
18211: waveform_sig_rx =350;
18212: waveform_sig_rx =607;
18213: waveform_sig_rx =381;
18214: waveform_sig_rx =547;
18215: waveform_sig_rx =398;
18216: waveform_sig_rx =592;
18217: waveform_sig_rx =276;
18218: waveform_sig_rx =598;
18219: waveform_sig_rx =489;
18220: waveform_sig_rx =227;
18221: waveform_sig_rx =693;
18222: waveform_sig_rx =337;
18223: waveform_sig_rx =270;
18224: waveform_sig_rx =651;
18225: waveform_sig_rx =309;
18226: waveform_sig_rx =269;
18227: waveform_sig_rx =589;
18228: waveform_sig_rx =337;
18229: waveform_sig_rx =279;
18230: waveform_sig_rx =431;
18231: waveform_sig_rx =460;
18232: waveform_sig_rx =225;
18233: waveform_sig_rx =322;
18234: waveform_sig_rx =525;
18235: waveform_sig_rx =199;
18236: waveform_sig_rx =229;
18237: waveform_sig_rx =469;
18238: waveform_sig_rx =293;
18239: waveform_sig_rx =144;
18240: waveform_sig_rx =476;
18241: waveform_sig_rx =278;
18242: waveform_sig_rx =161;
18243: waveform_sig_rx =337;
18244: waveform_sig_rx =370;
18245: waveform_sig_rx =169;
18246: waveform_sig_rx =162;
18247: waveform_sig_rx =407;
18248: waveform_sig_rx =185;
18249: waveform_sig_rx =89;
18250: waveform_sig_rx =416;
18251: waveform_sig_rx =200;
18252: waveform_sig_rx =86;
18253: waveform_sig_rx =319;
18254: waveform_sig_rx =85;
18255: waveform_sig_rx =274;
18256: waveform_sig_rx =124;
18257: waveform_sig_rx =263;
18258: waveform_sig_rx =-25;
18259: waveform_sig_rx =328;
18260: waveform_sig_rx =136;
18261: waveform_sig_rx =-36;
18262: waveform_sig_rx =377;
18263: waveform_sig_rx =-10;
18264: waveform_sig_rx =34;
18265: waveform_sig_rx =314;
18266: waveform_sig_rx =31;
18267: waveform_sig_rx =-21;
18268: waveform_sig_rx =234;
18269: waveform_sig_rx =103;
18270: waveform_sig_rx =-55;
18271: waveform_sig_rx =145;
18272: waveform_sig_rx =192;
18273: waveform_sig_rx =-169;
18274: waveform_sig_rx =90;
18275: waveform_sig_rx =200;
18276: waveform_sig_rx =-120;
18277: waveform_sig_rx =28;
18278: waveform_sig_rx =123;
18279: waveform_sig_rx =-25;
18280: waveform_sig_rx =-135;
18281: waveform_sig_rx =119;
18282: waveform_sig_rx =7;
18283: waveform_sig_rx =-147;
18284: waveform_sig_rx =14;
18285: waveform_sig_rx =84;
18286: waveform_sig_rx =-174;
18287: waveform_sig_rx =-126;
18288: waveform_sig_rx =121;
18289: waveform_sig_rx =-169;
18290: waveform_sig_rx =-195;
18291: waveform_sig_rx =123;
18292: waveform_sig_rx =-144;
18293: waveform_sig_rx =-186;
18294: waveform_sig_rx =23;
18295: waveform_sig_rx =-229;
18296: waveform_sig_rx =8;
18297: waveform_sig_rx =-178;
18298: waveform_sig_rx =-55;
18299: waveform_sig_rx =-289;
18300: waveform_sig_rx =13;
18301: waveform_sig_rx =-194;
18302: waveform_sig_rx =-276;
18303: waveform_sig_rx =8;
18304: waveform_sig_rx =-259;
18305: waveform_sig_rx =-299;
18306: waveform_sig_rx =-28;
18307: waveform_sig_rx =-217;
18308: waveform_sig_rx =-420;
18309: waveform_sig_rx =-15;
18310: waveform_sig_rx =-245;
18311: waveform_sig_rx =-418;
18312: waveform_sig_rx =-97;
18313: waveform_sig_rx =-196;
18314: waveform_sig_rx =-456;
18315: waveform_sig_rx =-191;
18316: waveform_sig_rx =-182;
18317: waveform_sig_rx =-398;
18318: waveform_sig_rx =-311;
18319: waveform_sig_rx =-196;
18320: waveform_sig_rx =-322;
18321: waveform_sig_rx =-453;
18322: waveform_sig_rx =-181;
18323: waveform_sig_rx =-294;
18324: waveform_sig_rx =-464;
18325: waveform_sig_rx =-302;
18326: waveform_sig_rx =-188;
18327: waveform_sig_rx =-529;
18328: waveform_sig_rx =-419;
18329: waveform_sig_rx =-161;
18330: waveform_sig_rx =-527;
18331: waveform_sig_rx =-452;
18332: waveform_sig_rx =-195;
18333: waveform_sig_rx =-486;
18334: waveform_sig_rx =-430;
18335: waveform_sig_rx =-352;
18336: waveform_sig_rx =-532;
18337: waveform_sig_rx =-291;
18338: waveform_sig_rx =-546;
18339: waveform_sig_rx =-336;
18340: waveform_sig_rx =-592;
18341: waveform_sig_rx =-339;
18342: waveform_sig_rx =-467;
18343: waveform_sig_rx =-637;
18344: waveform_sig_rx =-309;
18345: waveform_sig_rx =-527;
18346: waveform_sig_rx =-673;
18347: waveform_sig_rx =-256;
18348: waveform_sig_rx =-580;
18349: waveform_sig_rx =-707;
18350: waveform_sig_rx =-251;
18351: waveform_sig_rx =-610;
18352: waveform_sig_rx =-658;
18353: waveform_sig_rx =-391;
18354: waveform_sig_rx =-528;
18355: waveform_sig_rx =-716;
18356: waveform_sig_rx =-491;
18357: waveform_sig_rx =-464;
18358: waveform_sig_rx =-684;
18359: waveform_sig_rx =-613;
18360: waveform_sig_rx =-459;
18361: waveform_sig_rx =-620;
18362: waveform_sig_rx =-727;
18363: waveform_sig_rx =-473;
18364: waveform_sig_rx =-567;
18365: waveform_sig_rx =-787;
18366: waveform_sig_rx =-573;
18367: waveform_sig_rx =-448;
18368: waveform_sig_rx =-853;
18369: waveform_sig_rx =-608;
18370: waveform_sig_rx =-485;
18371: waveform_sig_rx =-814;
18372: waveform_sig_rx =-663;
18373: waveform_sig_rx =-560;
18374: waveform_sig_rx =-684;
18375: waveform_sig_rx =-733;
18376: waveform_sig_rx =-662;
18377: waveform_sig_rx =-701;
18378: waveform_sig_rx =-645;
18379: waveform_sig_rx =-782;
18380: waveform_sig_rx =-579;
18381: waveform_sig_rx =-901;
18382: waveform_sig_rx =-525;
18383: waveform_sig_rx =-782;
18384: waveform_sig_rx =-874;
18385: waveform_sig_rx =-519;
18386: waveform_sig_rx =-851;
18387: waveform_sig_rx =-896;
18388: waveform_sig_rx =-535;
18389: waveform_sig_rx =-867;
18390: waveform_sig_rx =-941;
18391: waveform_sig_rx =-504;
18392: waveform_sig_rx =-903;
18393: waveform_sig_rx =-903;
18394: waveform_sig_rx =-615;
18395: waveform_sig_rx =-823;
18396: waveform_sig_rx =-935;
18397: waveform_sig_rx =-760;
18398: waveform_sig_rx =-734;
18399: waveform_sig_rx =-904;
18400: waveform_sig_rx =-916;
18401: waveform_sig_rx =-660;
18402: waveform_sig_rx =-866;
18403: waveform_sig_rx =-1006;
18404: waveform_sig_rx =-635;
18405: waveform_sig_rx =-871;
18406: waveform_sig_rx =-989;
18407: waveform_sig_rx =-738;
18408: waveform_sig_rx =-770;
18409: waveform_sig_rx =-1017;
18410: waveform_sig_rx =-831;
18411: waveform_sig_rx =-755;
18412: waveform_sig_rx =-982;
18413: waveform_sig_rx =-940;
18414: waveform_sig_rx =-738;
18415: waveform_sig_rx =-921;
18416: waveform_sig_rx =-991;
18417: waveform_sig_rx =-844;
18418: waveform_sig_rx =-953;
18419: waveform_sig_rx =-904;
18420: waveform_sig_rx =-956;
18421: waveform_sig_rx =-830;
18422: waveform_sig_rx =-1131;
18423: waveform_sig_rx =-714;
18424: waveform_sig_rx =-1055;
18425: waveform_sig_rx =-1081;
18426: waveform_sig_rx =-721;
18427: waveform_sig_rx =-1119;
18428: waveform_sig_rx =-1061;
18429: waveform_sig_rx =-724;
18430: waveform_sig_rx =-1111;
18431: waveform_sig_rx =-1091;
18432: waveform_sig_rx =-753;
18433: waveform_sig_rx =-1121;
18434: waveform_sig_rx =-1053;
18435: waveform_sig_rx =-902;
18436: waveform_sig_rx =-974;
18437: waveform_sig_rx =-1124;
18438: waveform_sig_rx =-975;
18439: waveform_sig_rx =-865;
18440: waveform_sig_rx =-1139;
18441: waveform_sig_rx =-1081;
18442: waveform_sig_rx =-812;
18443: waveform_sig_rx =-1121;
18444: waveform_sig_rx =-1124;
18445: waveform_sig_rx =-853;
18446: waveform_sig_rx =-1085;
18447: waveform_sig_rx =-1100;
18448: waveform_sig_rx =-970;
18449: waveform_sig_rx =-946;
18450: waveform_sig_rx =-1182;
18451: waveform_sig_rx =-1028;
18452: waveform_sig_rx =-891;
18453: waveform_sig_rx =-1182;
18454: waveform_sig_rx =-1125;
18455: waveform_sig_rx =-874;
18456: waveform_sig_rx =-1122;
18457: waveform_sig_rx =-1128;
18458: waveform_sig_rx =-1000;
18459: waveform_sig_rx =-1122;
18460: waveform_sig_rx =-1027;
18461: waveform_sig_rx =-1100;
18462: waveform_sig_rx =-1027;
18463: waveform_sig_rx =-1269;
18464: waveform_sig_rx =-862;
18465: waveform_sig_rx =-1249;
18466: waveform_sig_rx =-1155;
18467: waveform_sig_rx =-885;
18468: waveform_sig_rx =-1292;
18469: waveform_sig_rx =-1108;
18470: waveform_sig_rx =-935;
18471: waveform_sig_rx =-1209;
18472: waveform_sig_rx =-1187;
18473: waveform_sig_rx =-934;
18474: waveform_sig_rx =-1181;
18475: waveform_sig_rx =-1209;
18476: waveform_sig_rx =-999;
18477: waveform_sig_rx =-1055;
18478: waveform_sig_rx =-1316;
18479: waveform_sig_rx =-1014;
18480: waveform_sig_rx =-1019;
18481: waveform_sig_rx =-1278;
18482: waveform_sig_rx =-1133;
18483: waveform_sig_rx =-987;
18484: waveform_sig_rx =-1232;
18485: waveform_sig_rx =-1217;
18486: waveform_sig_rx =-984;
18487: waveform_sig_rx =-1178;
18488: waveform_sig_rx =-1250;
18489: waveform_sig_rx =-1058;
18490: waveform_sig_rx =-1049;
18491: waveform_sig_rx =-1300;
18492: waveform_sig_rx =-1137;
18493: waveform_sig_rx =-992;
18494: waveform_sig_rx =-1284;
18495: waveform_sig_rx =-1224;
18496: waveform_sig_rx =-931;
18497: waveform_sig_rx =-1257;
18498: waveform_sig_rx =-1179;
18499: waveform_sig_rx =-1070;
18500: waveform_sig_rx =-1257;
18501: waveform_sig_rx =-1053;
18502: waveform_sig_rx =-1194;
18503: waveform_sig_rx =-1134;
18504: waveform_sig_rx =-1296;
18505: waveform_sig_rx =-968;
18506: waveform_sig_rx =-1303;
18507: waveform_sig_rx =-1202;
18508: waveform_sig_rx =-1016;
18509: waveform_sig_rx =-1298;
18510: waveform_sig_rx =-1216;
18511: waveform_sig_rx =-982;
18512: waveform_sig_rx =-1279;
18513: waveform_sig_rx =-1274;
18514: waveform_sig_rx =-930;
18515: waveform_sig_rx =-1271;
18516: waveform_sig_rx =-1258;
18517: waveform_sig_rx =-1027;
18518: waveform_sig_rx =-1139;
18519: waveform_sig_rx =-1358;
18520: waveform_sig_rx =-1032;
18521: waveform_sig_rx =-1084;
18522: waveform_sig_rx =-1310;
18523: waveform_sig_rx =-1152;
18524: waveform_sig_rx =-1035;
18525: waveform_sig_rx =-1255;
18526: waveform_sig_rx =-1202;
18527: waveform_sig_rx =-1028;
18528: waveform_sig_rx =-1164;
18529: waveform_sig_rx =-1282;
18530: waveform_sig_rx =-1085;
18531: waveform_sig_rx =-1027;
18532: waveform_sig_rx =-1372;
18533: waveform_sig_rx =-1103;
18534: waveform_sig_rx =-994;
18535: waveform_sig_rx =-1359;
18536: waveform_sig_rx =-1148;
18537: waveform_sig_rx =-985;
18538: waveform_sig_rx =-1301;
18539: waveform_sig_rx =-1110;
18540: waveform_sig_rx =-1159;
18541: waveform_sig_rx =-1208;
18542: waveform_sig_rx =-1065;
18543: waveform_sig_rx =-1218;
18544: waveform_sig_rx =-1058;
18545: waveform_sig_rx =-1292;
18546: waveform_sig_rx =-959;
18547: waveform_sig_rx =-1228;
18548: waveform_sig_rx =-1196;
18549: waveform_sig_rx =-934;
18550: waveform_sig_rx =-1270;
18551: waveform_sig_rx =-1187;
18552: waveform_sig_rx =-921;
18553: waveform_sig_rx =-1277;
18554: waveform_sig_rx =-1207;
18555: waveform_sig_rx =-894;
18556: waveform_sig_rx =-1246;
18557: waveform_sig_rx =-1199;
18558: waveform_sig_rx =-955;
18559: waveform_sig_rx =-1126;
18560: waveform_sig_rx =-1300;
18561: waveform_sig_rx =-929;
18562: waveform_sig_rx =-1097;
18563: waveform_sig_rx =-1211;
18564: waveform_sig_rx =-1099;
18565: waveform_sig_rx =-1005;
18566: waveform_sig_rx =-1146;
18567: waveform_sig_rx =-1195;
18568: waveform_sig_rx =-964;
18569: waveform_sig_rx =-1100;
18570: waveform_sig_rx =-1273;
18571: waveform_sig_rx =-931;
18572: waveform_sig_rx =-1029;
18573: waveform_sig_rx =-1300;
18574: waveform_sig_rx =-955;
18575: waveform_sig_rx =-988;
18576: waveform_sig_rx =-1224;
18577: waveform_sig_rx =-1060;
18578: waveform_sig_rx =-924;
18579: waveform_sig_rx =-1151;
18580: waveform_sig_rx =-1040;
18581: waveform_sig_rx =-1085;
18582: waveform_sig_rx =-1076;
18583: waveform_sig_rx =-1009;
18584: waveform_sig_rx =-1100;
18585: waveform_sig_rx =-966;
18586: waveform_sig_rx =-1216;
18587: waveform_sig_rx =-815;
18588: waveform_sig_rx =-1189;
18589: waveform_sig_rx =-1111;
18590: waveform_sig_rx =-820;
18591: waveform_sig_rx =-1204;
18592: waveform_sig_rx =-1070;
18593: waveform_sig_rx =-788;
18594: waveform_sig_rx =-1201;
18595: waveform_sig_rx =-1064;
18596: waveform_sig_rx =-770;
18597: waveform_sig_rx =-1172;
18598: waveform_sig_rx =-1045;
18599: waveform_sig_rx =-848;
18600: waveform_sig_rx =-1059;
18601: waveform_sig_rx =-1125;
18602: waveform_sig_rx =-840;
18603: waveform_sig_rx =-989;
18604: waveform_sig_rx =-1009;
18605: waveform_sig_rx =-1019;
18606: waveform_sig_rx =-823;
18607: waveform_sig_rx =-1027;
18608: waveform_sig_rx =-1091;
18609: waveform_sig_rx =-729;
18610: waveform_sig_rx =-1038;
18611: waveform_sig_rx =-1071;
18612: waveform_sig_rx =-766;
18613: waveform_sig_rx =-936;
18614: waveform_sig_rx =-1080;
18615: waveform_sig_rx =-852;
18616: waveform_sig_rx =-853;
18617: waveform_sig_rx =-1060;
18618: waveform_sig_rx =-943;
18619: waveform_sig_rx =-760;
18620: waveform_sig_rx =-1028;
18621: waveform_sig_rx =-890;
18622: waveform_sig_rx =-910;
18623: waveform_sig_rx =-907;
18624: waveform_sig_rx =-868;
18625: waveform_sig_rx =-914;
18626: waveform_sig_rx =-830;
18627: waveform_sig_rx =-1072;
18628: waveform_sig_rx =-626;
18629: waveform_sig_rx =-1058;
18630: waveform_sig_rx =-918;
18631: waveform_sig_rx =-626;
18632: waveform_sig_rx =-1111;
18633: waveform_sig_rx =-817;
18634: waveform_sig_rx =-636;
18635: waveform_sig_rx =-1067;
18636: waveform_sig_rx =-814;
18637: waveform_sig_rx =-657;
18638: waveform_sig_rx =-972;
18639: waveform_sig_rx =-830;
18640: waveform_sig_rx =-712;
18641: waveform_sig_rx =-805;
18642: waveform_sig_rx =-974;
18643: waveform_sig_rx =-646;
18644: waveform_sig_rx =-766;
18645: waveform_sig_rx =-899;
18646: waveform_sig_rx =-807;
18647: waveform_sig_rx =-591;
18648: waveform_sig_rx =-890;
18649: waveform_sig_rx =-852;
18650: waveform_sig_rx =-545;
18651: waveform_sig_rx =-891;
18652: waveform_sig_rx =-810;
18653: waveform_sig_rx =-588;
18654: waveform_sig_rx =-755;
18655: waveform_sig_rx =-818;
18656: waveform_sig_rx =-681;
18657: waveform_sig_rx =-611;
18658: waveform_sig_rx =-843;
18659: waveform_sig_rx =-755;
18660: waveform_sig_rx =-499;
18661: waveform_sig_rx =-847;
18662: waveform_sig_rx =-665;
18663: waveform_sig_rx =-692;
18664: waveform_sig_rx =-703;
18665: waveform_sig_rx =-626;
18666: waveform_sig_rx =-655;
18667: waveform_sig_rx =-644;
18668: waveform_sig_rx =-775;
18669: waveform_sig_rx =-391;
18670: waveform_sig_rx =-878;
18671: waveform_sig_rx =-611;
18672: waveform_sig_rx =-444;
18673: waveform_sig_rx =-886;
18674: waveform_sig_rx =-547;
18675: waveform_sig_rx =-478;
18676: waveform_sig_rx =-809;
18677: waveform_sig_rx =-558;
18678: waveform_sig_rx =-466;
18679: waveform_sig_rx =-697;
18680: waveform_sig_rx =-615;
18681: waveform_sig_rx =-463;
18682: waveform_sig_rx =-540;
18683: waveform_sig_rx =-758;
18684: waveform_sig_rx =-379;
18685: waveform_sig_rx =-515;
18686: waveform_sig_rx =-681;
18687: waveform_sig_rx =-507;
18688: waveform_sig_rx =-390;
18689: waveform_sig_rx =-679;
18690: waveform_sig_rx =-528;
18691: waveform_sig_rx =-357;
18692: waveform_sig_rx =-604;
18693: waveform_sig_rx =-557;
18694: waveform_sig_rx =-392;
18695: waveform_sig_rx =-468;
18696: waveform_sig_rx =-630;
18697: waveform_sig_rx =-432;
18698: waveform_sig_rx =-354;
18699: waveform_sig_rx =-639;
18700: waveform_sig_rx =-462;
18701: waveform_sig_rx =-249;
18702: waveform_sig_rx =-636;
18703: waveform_sig_rx =-368;
18704: waveform_sig_rx =-442;
18705: waveform_sig_rx =-456;
18706: waveform_sig_rx =-371;
18707: waveform_sig_rx =-413;
18708: waveform_sig_rx =-398;
18709: waveform_sig_rx =-500;
18710: waveform_sig_rx =-180;
18711: waveform_sig_rx =-616;
18712: waveform_sig_rx =-316;
18713: waveform_sig_rx =-244;
18714: waveform_sig_rx =-574;
18715: waveform_sig_rx =-275;
18716: waveform_sig_rx =-223;
18717: waveform_sig_rx =-485;
18718: waveform_sig_rx =-324;
18719: waveform_sig_rx =-161;
18720: waveform_sig_rx =-437;
18721: waveform_sig_rx =-366;
18722: waveform_sig_rx =-146;
18723: waveform_sig_rx =-307;
18724: waveform_sig_rx =-495;
18725: waveform_sig_rx =-52;
18726: waveform_sig_rx =-304;
18727: waveform_sig_rx =-380;
18728: waveform_sig_rx =-203;
18729: waveform_sig_rx =-170;
18730: waveform_sig_rx =-359;
18731: waveform_sig_rx =-252;
18732: waveform_sig_rx =-84;
18733: waveform_sig_rx =-277;
18734: waveform_sig_rx =-320;
18735: waveform_sig_rx =-66;
18736: waveform_sig_rx =-169;
18737: waveform_sig_rx =-373;
18738: waveform_sig_rx =-77;
18739: waveform_sig_rx =-82;
18740: waveform_sig_rx =-364;
18741: waveform_sig_rx =-141;
18742: waveform_sig_rx =-2;
18743: waveform_sig_rx =-334;
18744: waveform_sig_rx =-65;
18745: waveform_sig_rx =-167;
18746: waveform_sig_rx =-139;
18747: waveform_sig_rx =-76;
18748: waveform_sig_rx =-124;
18749: waveform_sig_rx =-128;
18750: waveform_sig_rx =-184;
18751: waveform_sig_rx =70;
18752: waveform_sig_rx =-281;
18753: waveform_sig_rx =-28;
18754: waveform_sig_rx =31;
18755: waveform_sig_rx =-215;
18756: waveform_sig_rx =-50;
18757: waveform_sig_rx =100;
18758: waveform_sig_rx =-234;
18759: waveform_sig_rx =-86;
18760: waveform_sig_rx =187;
18761: waveform_sig_rx =-236;
18762: waveform_sig_rx =-28;
18763: waveform_sig_rx =173;
18764: waveform_sig_rx =-109;
18765: waveform_sig_rx =-114;
18766: waveform_sig_rx =177;
18767: waveform_sig_rx =-24;
18768: waveform_sig_rx =-40;
18769: waveform_sig_rx =39;
18770: waveform_sig_rx =183;
18771: waveform_sig_rx =-70;
18772: waveform_sig_rx =40;
18773: waveform_sig_rx =226;
18774: waveform_sig_rx =-24;
18775: waveform_sig_rx =-21;
18776: waveform_sig_rx =240;
18777: waveform_sig_rx =125;
18778: waveform_sig_rx =-95;
18779: waveform_sig_rx =253;
18780: waveform_sig_rx =178;
18781: waveform_sig_rx =-61;
18782: waveform_sig_rx =226;
18783: waveform_sig_rx =254;
18784: waveform_sig_rx =-12;
18785: waveform_sig_rx =258;
18786: waveform_sig_rx =51;
18787: waveform_sig_rx =216;
18788: waveform_sig_rx =154;
18789: waveform_sig_rx =160;
18790: waveform_sig_rx =216;
18791: waveform_sig_rx =67;
18792: waveform_sig_rx =390;
18793: waveform_sig_rx =28;
18794: waveform_sig_rx =230;
18795: waveform_sig_rx =390;
18796: waveform_sig_rx =2;
18797: waveform_sig_rx =281;
18798: waveform_sig_rx =448;
18799: waveform_sig_rx =-12;
18800: waveform_sig_rx =301;
18801: waveform_sig_rx =457;
18802: waveform_sig_rx =57;
18803: waveform_sig_rx =322;
18804: waveform_sig_rx =407;
18805: waveform_sig_rx =200;
18806: waveform_sig_rx =175;
18807: waveform_sig_rx =452;
18808: waveform_sig_rx =286;
18809: waveform_sig_rx =220;
18810: waveform_sig_rx =337;
18811: waveform_sig_rx =455;
18812: waveform_sig_rx =188;
18813: waveform_sig_rx =327;
18814: waveform_sig_rx =517;
18815: waveform_sig_rx =262;
18816: waveform_sig_rx =234;
18817: waveform_sig_rx =570;
18818: waveform_sig_rx =356;
18819: waveform_sig_rx =198;
18820: waveform_sig_rx =574;
18821: waveform_sig_rx =386;
18822: waveform_sig_rx =276;
18823: waveform_sig_rx =459;
18824: waveform_sig_rx =498;
18825: waveform_sig_rx =334;
18826: waveform_sig_rx =448;
18827: waveform_sig_rx =392;
18828: waveform_sig_rx =508;
18829: waveform_sig_rx =371;
18830: waveform_sig_rx =531;
18831: waveform_sig_rx =438;
18832: waveform_sig_rx =371;
18833: waveform_sig_rx =718;
18834: waveform_sig_rx =227;
18835: waveform_sig_rx =566;
18836: waveform_sig_rx =647;
18837: waveform_sig_rx =240;
18838: waveform_sig_rx =621;
18839: waveform_sig_rx =652;
18840: waveform_sig_rx =277;
18841: waveform_sig_rx =593;
18842: waveform_sig_rx =709;
18843: waveform_sig_rx =333;
18844: waveform_sig_rx =597;
18845: waveform_sig_rx =675;
18846: waveform_sig_rx =468;
18847: waveform_sig_rx =469;
18848: waveform_sig_rx =715;
18849: waveform_sig_rx =570;
18850: waveform_sig_rx =481;
18851: waveform_sig_rx =592;
18852: waveform_sig_rx =770;
18853: waveform_sig_rx =412;
18854: waveform_sig_rx =610;
18855: waveform_sig_rx =799;
18856: waveform_sig_rx =451;
18857: waveform_sig_rx =583;
18858: waveform_sig_rx =820;
18859: waveform_sig_rx =560;
18860: waveform_sig_rx =544;
18861: waveform_sig_rx =779;
18862: waveform_sig_rx =672;
18863: waveform_sig_rx =574;
18864: waveform_sig_rx =678;
18865: waveform_sig_rx =835;
18866: waveform_sig_rx =547;
18867: waveform_sig_rx =697;
18868: waveform_sig_rx =676;
18869: waveform_sig_rx =693;
18870: waveform_sig_rx =679;
18871: waveform_sig_rx =808;
18872: waveform_sig_rx =629;
18873: waveform_sig_rx =703;
18874: waveform_sig_rx =923;
18875: waveform_sig_rx =466;
18876: waveform_sig_rx =883;
18877: waveform_sig_rx =832;
18878: waveform_sig_rx =523;
18879: waveform_sig_rx =890;
18880: waveform_sig_rx =885;
18881: waveform_sig_rx =504;
18882: waveform_sig_rx =888;
18883: waveform_sig_rx =893;
18884: waveform_sig_rx =582;
18885: waveform_sig_rx =891;
18886: waveform_sig_rx =832;
18887: waveform_sig_rx =772;
18888: waveform_sig_rx =672;
18889: waveform_sig_rx =935;
18890: waveform_sig_rx =859;
18891: waveform_sig_rx =635;
18892: waveform_sig_rx =898;
18893: waveform_sig_rx =973;
18894: waveform_sig_rx =590;
18895: waveform_sig_rx =931;
18896: waveform_sig_rx =936;
18897: waveform_sig_rx =723;
18898: waveform_sig_rx =826;
18899: waveform_sig_rx =980;
18900: waveform_sig_rx =857;
18901: waveform_sig_rx =716;
18902: waveform_sig_rx =1007;
18903: waveform_sig_rx =899;
18904: waveform_sig_rx =742;
18905: waveform_sig_rx =939;
18906: waveform_sig_rx =1040;
18907: waveform_sig_rx =737;
18908: waveform_sig_rx =972;
18909: waveform_sig_rx =898;
18910: waveform_sig_rx =886;
18911: waveform_sig_rx =908;
18912: waveform_sig_rx =983;
18913: waveform_sig_rx =806;
18914: waveform_sig_rx =944;
18915: waveform_sig_rx =1076;
18916: waveform_sig_rx =677;
18917: waveform_sig_rx =1114;
18918: waveform_sig_rx =992;
18919: waveform_sig_rx =757;
18920: waveform_sig_rx =1111;
18921: waveform_sig_rx =1030;
18922: waveform_sig_rx =780;
18923: waveform_sig_rx =1046;
18924: waveform_sig_rx =1088;
18925: waveform_sig_rx =812;
18926: waveform_sig_rx =1001;
18927: waveform_sig_rx =1091;
18928: waveform_sig_rx =935;
18929: waveform_sig_rx =830;
18930: waveform_sig_rx =1192;
18931: waveform_sig_rx =945;
18932: waveform_sig_rx =840;
18933: waveform_sig_rx =1111;
18934: waveform_sig_rx =1053;
18935: waveform_sig_rx =835;
18936: waveform_sig_rx =1092;
18937: waveform_sig_rx =1059;
18938: waveform_sig_rx =937;
18939: waveform_sig_rx =951;
18940: waveform_sig_rx =1155;
18941: waveform_sig_rx =1018;
18942: waveform_sig_rx =846;
18943: waveform_sig_rx =1201;
18944: waveform_sig_rx =1050;
18945: waveform_sig_rx =852;
18946: waveform_sig_rx =1135;
18947: waveform_sig_rx =1152;
18948: waveform_sig_rx =865;
18949: waveform_sig_rx =1172;
18950: waveform_sig_rx =991;
18951: waveform_sig_rx =1053;
18952: waveform_sig_rx =1083;
18953: waveform_sig_rx =1081;
18954: waveform_sig_rx =973;
18955: waveform_sig_rx =1099;
18956: waveform_sig_rx =1166;
18957: waveform_sig_rx =867;
18958: waveform_sig_rx =1213;
18959: waveform_sig_rx =1094;
18960: waveform_sig_rx =938;
18961: waveform_sig_rx =1184;
18962: waveform_sig_rx =1195;
18963: waveform_sig_rx =873;
18964: waveform_sig_rx =1157;
18965: waveform_sig_rx =1247;
18966: waveform_sig_rx =887;
18967: waveform_sig_rx =1148;
18968: waveform_sig_rx =1242;
18969: waveform_sig_rx =983;
18970: waveform_sig_rx =1003;
18971: waveform_sig_rx =1310;
18972: waveform_sig_rx =999;
18973: waveform_sig_rx =1019;
18974: waveform_sig_rx =1202;
18975: waveform_sig_rx =1162;
18976: waveform_sig_rx =971;
18977: waveform_sig_rx =1169;
18978: waveform_sig_rx =1204;
18979: waveform_sig_rx =1031;
18980: waveform_sig_rx =1043;
18981: waveform_sig_rx =1294;
18982: waveform_sig_rx =1083;
18983: waveform_sig_rx =937;
18984: waveform_sig_rx =1334;
18985: waveform_sig_rx =1110;
18986: waveform_sig_rx =960;
18987: waveform_sig_rx =1274;
18988: waveform_sig_rx =1189;
18989: waveform_sig_rx =981;
18990: waveform_sig_rx =1268;
18991: waveform_sig_rx =997;
18992: waveform_sig_rx =1229;
18993: waveform_sig_rx =1094;
18994: waveform_sig_rx =1164;
18995: waveform_sig_rx =1092;
18996: waveform_sig_rx =1126;
18997: waveform_sig_rx =1275;
18998: waveform_sig_rx =925;
18999: waveform_sig_rx =1262;
19000: waveform_sig_rx =1218;
19001: waveform_sig_rx =951;
19002: waveform_sig_rx =1264;
19003: waveform_sig_rx =1246;
19004: waveform_sig_rx =896;
19005: waveform_sig_rx =1259;
19006: waveform_sig_rx =1268;
19007: waveform_sig_rx =926;
19008: waveform_sig_rx =1213;
19009: waveform_sig_rx =1288;
19010: waveform_sig_rx =994;
19011: waveform_sig_rx =1121;
19012: waveform_sig_rx =1341;
19013: waveform_sig_rx =1047;
19014: waveform_sig_rx =1129;
19015: waveform_sig_rx =1179;
19016: waveform_sig_rx =1244;
19017: waveform_sig_rx =1003;
19018: waveform_sig_rx =1164;
19019: waveform_sig_rx =1308;
19020: waveform_sig_rx =981;
19021: waveform_sig_rx =1085;
19022: waveform_sig_rx =1353;
19023: waveform_sig_rx =1001;
19024: waveform_sig_rx =1024;
19025: waveform_sig_rx =1340;
19026: waveform_sig_rx =1067;
19027: waveform_sig_rx =1024;
19028: waveform_sig_rx =1256;
19029: waveform_sig_rx =1201;
19030: waveform_sig_rx =1014;
19031: waveform_sig_rx =1232;
19032: waveform_sig_rx =1040;
19033: waveform_sig_rx =1266;
19034: waveform_sig_rx =1074;
19035: waveform_sig_rx =1235;
19036: waveform_sig_rx =1063;
19037: waveform_sig_rx =1133;
19038: waveform_sig_rx =1312;
19039: waveform_sig_rx =876;
19040: waveform_sig_rx =1274;
19041: waveform_sig_rx =1217;
19042: waveform_sig_rx =883;
19043: waveform_sig_rx =1321;
19044: waveform_sig_rx =1198;
19045: waveform_sig_rx =861;
19046: waveform_sig_rx =1299;
19047: waveform_sig_rx =1183;
19048: waveform_sig_rx =902;
19049: waveform_sig_rx =1222;
19050: waveform_sig_rx =1178;
19051: waveform_sig_rx =969;
19052: waveform_sig_rx =1091;
19053: waveform_sig_rx =1243;
19054: waveform_sig_rx =1043;
19055: waveform_sig_rx =1039;
19056: waveform_sig_rx =1136;
19057: waveform_sig_rx =1243;
19058: waveform_sig_rx =907;
19059: waveform_sig_rx =1196;
19060: waveform_sig_rx =1260;
19061: waveform_sig_rx =911;
19062: waveform_sig_rx =1131;
19063: waveform_sig_rx =1275;
19064: waveform_sig_rx =965;
19065: waveform_sig_rx =1044;
19066: waveform_sig_rx =1224;
19067: waveform_sig_rx =1062;
19068: waveform_sig_rx =975;
19069: waveform_sig_rx =1176;
19070: waveform_sig_rx =1148;
19071: waveform_sig_rx =938;
19072: waveform_sig_rx =1157;
19073: waveform_sig_rx =995;
19074: waveform_sig_rx =1148;
19075: waveform_sig_rx =979;
19076: waveform_sig_rx =1190;
19077: waveform_sig_rx =926;
19078: waveform_sig_rx =1077;
19079: waveform_sig_rx =1202;
19080: waveform_sig_rx =776;
19081: waveform_sig_rx =1258;
19082: waveform_sig_rx =1081;
19083: waveform_sig_rx =797;
19084: waveform_sig_rx =1302;
19085: waveform_sig_rx =1026;
19086: waveform_sig_rx =833;
19087: waveform_sig_rx =1239;
19088: waveform_sig_rx =1038;
19089: waveform_sig_rx =888;
19090: waveform_sig_rx =1122;
19091: waveform_sig_rx =1096;
19092: waveform_sig_rx =924;
19093: waveform_sig_rx =956;
19094: waveform_sig_rx =1179;
19095: waveform_sig_rx =946;
19096: waveform_sig_rx =907;
19097: waveform_sig_rx =1095;
19098: waveform_sig_rx =1107;
19099: waveform_sig_rx =787;
19100: waveform_sig_rx =1119;
19101: waveform_sig_rx =1082;
19102: waveform_sig_rx =793;
19103: waveform_sig_rx =1038;
19104: waveform_sig_rx =1094;
19105: waveform_sig_rx =881;
19106: waveform_sig_rx =909;
19107: waveform_sig_rx =1080;
19108: waveform_sig_rx =975;
19109: waveform_sig_rx =797;
19110: waveform_sig_rx =1045;
19111: waveform_sig_rx =1041;
19112: waveform_sig_rx =755;
19113: waveform_sig_rx =1054;
19114: waveform_sig_rx =850;
19115: waveform_sig_rx =982;
19116: waveform_sig_rx =889;
19117: waveform_sig_rx =1022;
19118: waveform_sig_rx =739;
19119: waveform_sig_rx =1030;
19120: waveform_sig_rx =972;
19121: waveform_sig_rx =651;
19122: waveform_sig_rx =1146;
19123: waveform_sig_rx =825;
19124: waveform_sig_rx =728;
19125: waveform_sig_rx =1110;
19126: waveform_sig_rx =846;
19127: waveform_sig_rx =737;
19128: waveform_sig_rx =1014;
19129: waveform_sig_rx =894;
19130: waveform_sig_rx =762;
19131: waveform_sig_rx =913;
19132: waveform_sig_rx =990;
19133: waveform_sig_rx =735;
19134: waveform_sig_rx =792;
19135: waveform_sig_rx =1036;
19136: waveform_sig_rx =735;
19137: waveform_sig_rx =751;
19138: waveform_sig_rx =935;
19139: waveform_sig_rx =861;
19140: waveform_sig_rx =623;
19141: waveform_sig_rx =961;
19142: waveform_sig_rx =823;
19143: waveform_sig_rx =664;
19144: waveform_sig_rx =842;
19145: waveform_sig_rx =858;
19146: waveform_sig_rx =732;
19147: waveform_sig_rx =660;
19148: waveform_sig_rx =912;
19149: waveform_sig_rx =779;
19150: waveform_sig_rx =561;
19151: waveform_sig_rx =958;
19152: waveform_sig_rx =782;
19153: waveform_sig_rx =560;
19154: waveform_sig_rx =909;
19155: waveform_sig_rx =589;
19156: waveform_sig_rx =834;
19157: waveform_sig_rx =675;
19158: waveform_sig_rx =795;
19159: waveform_sig_rx =568;
19160: waveform_sig_rx =817;
19161: waveform_sig_rx =743;
19162: waveform_sig_rx =500;
19163: waveform_sig_rx =913;
19164: waveform_sig_rx =620;
19165: waveform_sig_rx =552;
19166: waveform_sig_rx =867;
19167: waveform_sig_rx =632;
19168: waveform_sig_rx =512;
19169: waveform_sig_rx =757;
19170: waveform_sig_rx =693;
19171: waveform_sig_rx =488;
19172: waveform_sig_rx =676;
19173: waveform_sig_rx =778;
19174: waveform_sig_rx =421;
19175: waveform_sig_rx =611;
19176: waveform_sig_rx =815;
19177: waveform_sig_rx =442;
19178: waveform_sig_rx =583;
19179: waveform_sig_rx =670;
19180: waveform_sig_rx =600;
19181: waveform_sig_rx =431;
19182: waveform_sig_rx =665;
19183: waveform_sig_rx =630;
19184: waveform_sig_rx =427;
19185: waveform_sig_rx =558;
19186: waveform_sig_rx =680;
19187: waveform_sig_rx =449;
19188: waveform_sig_rx =427;
19189: waveform_sig_rx =717;
19190: waveform_sig_rx =470;
19191: waveform_sig_rx =341;
19192: waveform_sig_rx =694;
19193: waveform_sig_rx =476;
19194: waveform_sig_rx =354;
19195: waveform_sig_rx =649;
19196: waveform_sig_rx =313;
19197: waveform_sig_rx =594;
19198: waveform_sig_rx =404;
19199: waveform_sig_rx =529;
19200: waveform_sig_rx =335;
19201: waveform_sig_rx =544;
19202: waveform_sig_rx =469;
19203: waveform_sig_rx =279;
19204: waveform_sig_rx =594;
19205: waveform_sig_rx =359;
19206: waveform_sig_rx =290;
19207: waveform_sig_rx =561;
19208: waveform_sig_rx =436;
19209: waveform_sig_rx =201;
19210: waveform_sig_rx =540;
19211: waveform_sig_rx =462;
19212: waveform_sig_rx =166;
19213: waveform_sig_rx =519;
19214: waveform_sig_rx =469;
19215: waveform_sig_rx =151;
19216: waveform_sig_rx =410;
19217: waveform_sig_rx =456;
19218: waveform_sig_rx =229;
19219: waveform_sig_rx =321;
19220: waveform_sig_rx =385;
19221: waveform_sig_rx =364;
19222: waveform_sig_rx =115;
19223: waveform_sig_rx =403;
19224: waveform_sig_rx =346;
19225: waveform_sig_rx =115;
19226: waveform_sig_rx =282;
19227: waveform_sig_rx =409;
19228: waveform_sig_rx =137;
19229: waveform_sig_rx =172;
19230: waveform_sig_rx =450;
19231: waveform_sig_rx =133;
19232: waveform_sig_rx =110;
19233: waveform_sig_rx =411;
19234: waveform_sig_rx =143;
19235: waveform_sig_rx =131;
19236: waveform_sig_rx =312;
19237: waveform_sig_rx =46;
19238: waveform_sig_rx =352;
19239: waveform_sig_rx =67;
19240: waveform_sig_rx =293;
19241: waveform_sig_rx =41;
19242: waveform_sig_rx =238;
19243: waveform_sig_rx =232;
19244: waveform_sig_rx =-46;
19245: waveform_sig_rx =304;
19246: waveform_sig_rx =152;
19247: waveform_sig_rx =-85;
19248: waveform_sig_rx =357;
19249: waveform_sig_rx =86;
19250: waveform_sig_rx =-136;
19251: waveform_sig_rx =358;
19252: waveform_sig_rx =45;
19253: waveform_sig_rx =-103;
19254: waveform_sig_rx =202;
19255: waveform_sig_rx =80;
19256: waveform_sig_rx =-109;
19257: waveform_sig_rx =83;
19258: waveform_sig_rx =157;
19259: waveform_sig_rx =-57;
19260: waveform_sig_rx =-33;
19261: waveform_sig_rx =125;
19262: waveform_sig_rx =45;
19263: waveform_sig_rx =-168;
19264: waveform_sig_rx =123;
19265: waveform_sig_rx =41;
19266: waveform_sig_rx =-200;
19267: waveform_sig_rx =3;
19268: waveform_sig_rx =150;
19269: waveform_sig_rx =-234;
19270: waveform_sig_rx =-49;
19271: waveform_sig_rx =113;
19272: waveform_sig_rx =-214;
19273: waveform_sig_rx =-94;
19274: waveform_sig_rx =3;
19275: waveform_sig_rx =-76;
19276: waveform_sig_rx =-154;
19277: waveform_sig_rx =-87;
19278: waveform_sig_rx =-131;
19279: waveform_sig_rx =-60;
19280: waveform_sig_rx =-216;
19281: waveform_sig_rx =13;
19282: waveform_sig_rx =-343;
19283: waveform_sig_rx =-2;
19284: waveform_sig_rx =-137;
19285: waveform_sig_rx =-403;
19286: waveform_sig_rx =62;
19287: waveform_sig_rx =-276;
19288: waveform_sig_rx =-345;
19289: waveform_sig_rx =35;
19290: waveform_sig_rx =-290;
19291: waveform_sig_rx =-403;
19292: waveform_sig_rx =12;
19293: waveform_sig_rx =-279;
19294: waveform_sig_rx =-384;
19295: waveform_sig_rx =-97;
19296: waveform_sig_rx =-224;
19297: waveform_sig_rx =-398;
19298: waveform_sig_rx =-239;
19299: waveform_sig_rx =-181;
19300: waveform_sig_rx =-355;
19301: waveform_sig_rx =-362;
19302: waveform_sig_rx =-179;
19303: waveform_sig_rx =-266;
19304: waveform_sig_rx =-504;
19305: waveform_sig_rx =-134;
19306: waveform_sig_rx =-285;
19307: waveform_sig_rx =-526;
19308: waveform_sig_rx =-216;
19309: waveform_sig_rx =-252;
19310: waveform_sig_rx =-509;
19311: waveform_sig_rx =-336;
19312: waveform_sig_rx =-246;
19313: waveform_sig_rx =-428;
19314: waveform_sig_rx =-465;
19315: waveform_sig_rx =-282;
19316: waveform_sig_rx =-328;
19317: waveform_sig_rx =-544;
19318: waveform_sig_rx =-300;
19319: waveform_sig_rx =-452;
19320: waveform_sig_rx =-393;
19321: waveform_sig_rx =-440;
19322: waveform_sig_rx =-345;
19323: waveform_sig_rx =-634;
19324: waveform_sig_rx =-244;
19325: waveform_sig_rx =-506;
19326: waveform_sig_rx =-610;
19327: waveform_sig_rx =-254;
19328: waveform_sig_rx =-600;
19329: waveform_sig_rx =-606;
19330: waveform_sig_rx =-264;
19331: waveform_sig_rx =-560;
19332: waveform_sig_rx =-706;
19333: waveform_sig_rx =-278;
19334: waveform_sig_rx =-601;
19335: waveform_sig_rx =-635;
19336: waveform_sig_rx =-405;
19337: waveform_sig_rx =-519;
19338: waveform_sig_rx =-666;
19339: waveform_sig_rx =-585;
19340: waveform_sig_rx =-418;
19341: waveform_sig_rx =-661;
19342: waveform_sig_rx =-688;
19343: waveform_sig_rx =-369;
19344: waveform_sig_rx =-648;
19345: waveform_sig_rx =-739;
19346: waveform_sig_rx =-383;
19347: waveform_sig_rx =-654;
19348: waveform_sig_rx =-703;
19349: waveform_sig_rx =-558;
19350: waveform_sig_rx =-518;
19351: waveform_sig_rx =-724;
19352: waveform_sig_rx =-706;
19353: waveform_sig_rx =-460;
19354: waveform_sig_rx =-724;
19355: waveform_sig_rx =-772;
19356: waveform_sig_rx =-482;
19357: waveform_sig_rx =-691;
19358: waveform_sig_rx =-789;
19359: waveform_sig_rx =-570;
19360: waveform_sig_rx =-788;
19361: waveform_sig_rx =-627;
19362: waveform_sig_rx =-730;
19363: waveform_sig_rx =-655;
19364: waveform_sig_rx =-879;
19365: waveform_sig_rx =-520;
19366: waveform_sig_rx =-797;
19367: waveform_sig_rx =-845;
19368: waveform_sig_rx =-528;
19369: waveform_sig_rx =-874;
19370: waveform_sig_rx =-826;
19371: waveform_sig_rx =-556;
19372: waveform_sig_rx =-846;
19373: waveform_sig_rx =-898;
19374: waveform_sig_rx =-578;
19375: waveform_sig_rx =-822;
19376: waveform_sig_rx =-895;
19377: waveform_sig_rx =-695;
19378: waveform_sig_rx =-676;
19379: waveform_sig_rx =-979;
19380: waveform_sig_rx =-779;
19381: waveform_sig_rx =-628;
19382: waveform_sig_rx =-981;
19383: waveform_sig_rx =-827;
19384: waveform_sig_rx =-648;
19385: waveform_sig_rx =-905;
19386: waveform_sig_rx =-903;
19387: waveform_sig_rx =-700;
19388: waveform_sig_rx =-818;
19389: waveform_sig_rx =-938;
19390: waveform_sig_rx =-832;
19391: waveform_sig_rx =-690;
19392: waveform_sig_rx =-1030;
19393: waveform_sig_rx =-905;
19394: waveform_sig_rx =-677;
19395: waveform_sig_rx =-1010;
19396: waveform_sig_rx =-957;
19397: waveform_sig_rx =-686;
19398: waveform_sig_rx =-950;
19399: waveform_sig_rx =-964;
19400: waveform_sig_rx =-799;
19401: waveform_sig_rx =-1009;
19402: waveform_sig_rx =-815;
19403: waveform_sig_rx =-953;
19404: waveform_sig_rx =-886;
19405: waveform_sig_rx =-1063;
19406: waveform_sig_rx =-746;
19407: waveform_sig_rx =-1037;
19408: waveform_sig_rx =-1021;
19409: waveform_sig_rx =-782;
19410: waveform_sig_rx =-1039;
19411: waveform_sig_rx =-1013;
19412: waveform_sig_rx =-775;
19413: waveform_sig_rx =-999;
19414: waveform_sig_rx =-1128;
19415: waveform_sig_rx =-746;
19416: waveform_sig_rx =-1010;
19417: waveform_sig_rx =-1139;
19418: waveform_sig_rx =-831;
19419: waveform_sig_rx =-927;
19420: waveform_sig_rx =-1214;
19421: waveform_sig_rx =-897;
19422: waveform_sig_rx =-886;
19423: waveform_sig_rx =-1155;
19424: waveform_sig_rx =-1010;
19425: waveform_sig_rx =-909;
19426: waveform_sig_rx =-1054;
19427: waveform_sig_rx =-1106;
19428: waveform_sig_rx =-924;
19429: waveform_sig_rx =-996;
19430: waveform_sig_rx =-1163;
19431: waveform_sig_rx =-988;
19432: waveform_sig_rx =-860;
19433: waveform_sig_rx =-1255;
19434: waveform_sig_rx =-1031;
19435: waveform_sig_rx =-877;
19436: waveform_sig_rx =-1214;
19437: waveform_sig_rx =-1077;
19438: waveform_sig_rx =-890;
19439: waveform_sig_rx =-1148;
19440: waveform_sig_rx =-1102;
19441: waveform_sig_rx =-1005;
19442: waveform_sig_rx =-1158;
19443: waveform_sig_rx =-961;
19444: waveform_sig_rx =-1161;
19445: waveform_sig_rx =-1015;
19446: waveform_sig_rx =-1207;
19447: waveform_sig_rx =-926;
19448: waveform_sig_rx =-1141;
19449: waveform_sig_rx =-1181;
19450: waveform_sig_rx =-938;
19451: waveform_sig_rx =-1160;
19452: waveform_sig_rx =-1222;
19453: waveform_sig_rx =-881;
19454: waveform_sig_rx =-1179;
19455: waveform_sig_rx =-1307;
19456: waveform_sig_rx =-802;
19457: waveform_sig_rx =-1207;
19458: waveform_sig_rx =-1231;
19459: waveform_sig_rx =-910;
19460: waveform_sig_rx =-1140;
19461: waveform_sig_rx =-1266;
19462: waveform_sig_rx =-1001;
19463: waveform_sig_rx =-1065;
19464: waveform_sig_rx =-1197;
19465: waveform_sig_rx =-1138;
19466: waveform_sig_rx =-1002;
19467: waveform_sig_rx =-1135;
19468: waveform_sig_rx =-1251;
19469: waveform_sig_rx =-970;
19470: waveform_sig_rx =-1108;
19471: waveform_sig_rx =-1322;
19472: waveform_sig_rx =-1012;
19473: waveform_sig_rx =-1031;
19474: waveform_sig_rx =-1360;
19475: waveform_sig_rx =-1051;
19476: waveform_sig_rx =-1015;
19477: waveform_sig_rx =-1297;
19478: waveform_sig_rx =-1152;
19479: waveform_sig_rx =-996;
19480: waveform_sig_rx =-1214;
19481: waveform_sig_rx =-1176;
19482: waveform_sig_rx =-1119;
19483: waveform_sig_rx =-1193;
19484: waveform_sig_rx =-1090;
19485: waveform_sig_rx =-1229;
19486: waveform_sig_rx =-1031;
19487: waveform_sig_rx =-1335;
19488: waveform_sig_rx =-963;
19489: waveform_sig_rx =-1219;
19490: waveform_sig_rx =-1305;
19491: waveform_sig_rx =-944;
19492: waveform_sig_rx =-1282;
19493: waveform_sig_rx =-1269;
19494: waveform_sig_rx =-873;
19495: waveform_sig_rx =-1304;
19496: waveform_sig_rx =-1291;
19497: waveform_sig_rx =-877;
19498: waveform_sig_rx =-1335;
19499: waveform_sig_rx =-1217;
19500: waveform_sig_rx =-1012;
19501: waveform_sig_rx =-1193;
19502: waveform_sig_rx =-1277;
19503: waveform_sig_rx =-1076;
19504: waveform_sig_rx =-1085;
19505: waveform_sig_rx =-1224;
19506: waveform_sig_rx =-1224;
19507: waveform_sig_rx =-979;
19508: waveform_sig_rx =-1200;
19509: waveform_sig_rx =-1308;
19510: waveform_sig_rx =-947;
19511: waveform_sig_rx =-1200;
19512: waveform_sig_rx =-1307;
19513: waveform_sig_rx =-1006;
19514: waveform_sig_rx =-1098;
19515: waveform_sig_rx =-1310;
19516: waveform_sig_rx =-1078;
19517: waveform_sig_rx =-1046;
19518: waveform_sig_rx =-1265;
19519: waveform_sig_rx =-1189;
19520: waveform_sig_rx =-1002;
19521: waveform_sig_rx =-1212;
19522: waveform_sig_rx =-1174;
19523: waveform_sig_rx =-1121;
19524: waveform_sig_rx =-1153;
19525: waveform_sig_rx =-1108;
19526: waveform_sig_rx =-1173;
19527: waveform_sig_rx =-1029;
19528: waveform_sig_rx =-1363;
19529: waveform_sig_rx =-884;
19530: waveform_sig_rx =-1256;
19531: waveform_sig_rx =-1239;
19532: waveform_sig_rx =-864;
19533: waveform_sig_rx =-1353;
19534: waveform_sig_rx =-1142;
19535: waveform_sig_rx =-889;
19536: waveform_sig_rx =-1318;
19537: waveform_sig_rx =-1139;
19538: waveform_sig_rx =-935;
19539: waveform_sig_rx =-1236;
19540: waveform_sig_rx =-1162;
19541: waveform_sig_rx =-1010;
19542: waveform_sig_rx =-1059;
19543: waveform_sig_rx =-1292;
19544: waveform_sig_rx =-993;
19545: waveform_sig_rx =-1030;
19546: waveform_sig_rx =-1225;
19547: waveform_sig_rx =-1134;
19548: waveform_sig_rx =-932;
19549: waveform_sig_rx =-1179;
19550: waveform_sig_rx =-1236;
19551: waveform_sig_rx =-884;
19552: waveform_sig_rx =-1166;
19553: waveform_sig_rx =-1227;
19554: waveform_sig_rx =-940;
19555: waveform_sig_rx =-1071;
19556: waveform_sig_rx =-1192;
19557: waveform_sig_rx =-1042;
19558: waveform_sig_rx =-986;
19559: waveform_sig_rx =-1151;
19560: waveform_sig_rx =-1160;
19561: waveform_sig_rx =-863;
19562: waveform_sig_rx =-1166;
19563: waveform_sig_rx =-1123;
19564: waveform_sig_rx =-981;
19565: waveform_sig_rx =-1137;
19566: waveform_sig_rx =-1013;
19567: waveform_sig_rx =-1065;
19568: waveform_sig_rx =-1009;
19569: waveform_sig_rx =-1212;
19570: waveform_sig_rx =-795;
19571: waveform_sig_rx =-1235;
19572: waveform_sig_rx =-1047;
19573: waveform_sig_rx =-819;
19574: waveform_sig_rx =-1247;
19575: waveform_sig_rx =-977;
19576: waveform_sig_rx =-873;
19577: waveform_sig_rx =-1166;
19578: waveform_sig_rx =-1051;
19579: waveform_sig_rx =-844;
19580: waveform_sig_rx =-1095;
19581: waveform_sig_rx =-1068;
19582: waveform_sig_rx =-876;
19583: waveform_sig_rx =-964;
19584: waveform_sig_rx =-1187;
19585: waveform_sig_rx =-850;
19586: waveform_sig_rx =-922;
19587: waveform_sig_rx =-1095;
19588: waveform_sig_rx =-991;
19589: waveform_sig_rx =-801;
19590: waveform_sig_rx =-1090;
19591: waveform_sig_rx =-1041;
19592: waveform_sig_rx =-766;
19593: waveform_sig_rx =-1055;
19594: waveform_sig_rx =-1014;
19595: waveform_sig_rx =-846;
19596: waveform_sig_rx =-896;
19597: waveform_sig_rx =-1044;
19598: waveform_sig_rx =-952;
19599: waveform_sig_rx =-750;
19600: waveform_sig_rx =-1074;
19601: waveform_sig_rx =-988;
19602: waveform_sig_rx =-662;
19603: waveform_sig_rx =-1108;
19604: waveform_sig_rx =-858;
19605: waveform_sig_rx =-865;
19606: waveform_sig_rx =-1001;
19607: waveform_sig_rx =-780;
19608: waveform_sig_rx =-918;
19609: waveform_sig_rx =-846;
19610: waveform_sig_rx =-986;
19611: waveform_sig_rx =-650;
19612: waveform_sig_rx =-1013;
19613: waveform_sig_rx =-867;
19614: waveform_sig_rx =-666;
19615: waveform_sig_rx =-1040;
19616: waveform_sig_rx =-819;
19617: waveform_sig_rx =-658;
19618: waveform_sig_rx =-995;
19619: waveform_sig_rx =-872;
19620: waveform_sig_rx =-656;
19621: waveform_sig_rx =-925;
19622: waveform_sig_rx =-900;
19623: waveform_sig_rx =-675;
19624: waveform_sig_rx =-779;
19625: waveform_sig_rx =-1020;
19626: waveform_sig_rx =-598;
19627: waveform_sig_rx =-765;
19628: waveform_sig_rx =-917;
19629: waveform_sig_rx =-727;
19630: waveform_sig_rx =-664;
19631: waveform_sig_rx =-848;
19632: waveform_sig_rx =-808;
19633: waveform_sig_rx =-621;
19634: waveform_sig_rx =-784;
19635: waveform_sig_rx =-869;
19636: waveform_sig_rx =-638;
19637: waveform_sig_rx =-653;
19638: waveform_sig_rx =-932;
19639: waveform_sig_rx =-642;
19640: waveform_sig_rx =-577;
19641: waveform_sig_rx =-924;
19642: waveform_sig_rx =-688;
19643: waveform_sig_rx =-531;
19644: waveform_sig_rx =-872;
19645: waveform_sig_rx =-633;
19646: waveform_sig_rx =-685;
19647: waveform_sig_rx =-716;
19648: waveform_sig_rx =-600;
19649: waveform_sig_rx =-711;
19650: waveform_sig_rx =-597;
19651: waveform_sig_rx =-779;
19652: waveform_sig_rx =-442;
19653: waveform_sig_rx =-803;
19654: waveform_sig_rx =-656;
19655: waveform_sig_rx =-475;
19656: waveform_sig_rx =-795;
19657: waveform_sig_rx =-623;
19658: waveform_sig_rx =-445;
19659: waveform_sig_rx =-757;
19660: waveform_sig_rx =-678;
19661: waveform_sig_rx =-352;
19662: waveform_sig_rx =-732;
19663: waveform_sig_rx =-657;
19664: waveform_sig_rx =-366;
19665: waveform_sig_rx =-628;
19666: waveform_sig_rx =-717;
19667: waveform_sig_rx =-360;
19668: waveform_sig_rx =-601;
19669: waveform_sig_rx =-596;
19670: waveform_sig_rx =-541;
19671: waveform_sig_rx =-422;
19672: waveform_sig_rx =-568;
19673: waveform_sig_rx =-622;
19674: waveform_sig_rx =-306;
19675: waveform_sig_rx =-565;
19676: waveform_sig_rx =-640;
19677: waveform_sig_rx =-311;
19678: waveform_sig_rx =-461;
19679: waveform_sig_rx =-647;
19680: waveform_sig_rx =-362;
19681: waveform_sig_rx =-365;
19682: waveform_sig_rx =-618;
19683: waveform_sig_rx =-411;
19684: waveform_sig_rx =-298;
19685: waveform_sig_rx =-584;
19686: waveform_sig_rx =-370;
19687: waveform_sig_rx =-483;
19688: waveform_sig_rx =-402;
19689: waveform_sig_rx =-369;
19690: waveform_sig_rx =-459;
19691: waveform_sig_rx =-315;
19692: waveform_sig_rx =-562;
19693: waveform_sig_rx =-161;
19694: waveform_sig_rx =-521;
19695: waveform_sig_rx =-409;
19696: waveform_sig_rx =-152;
19697: waveform_sig_rx =-536;
19698: waveform_sig_rx =-351;
19699: waveform_sig_rx =-109;
19700: waveform_sig_rx =-535;
19701: waveform_sig_rx =-328;
19702: waveform_sig_rx =-78;
19703: waveform_sig_rx =-530;
19704: waveform_sig_rx =-290;
19705: waveform_sig_rx =-146;
19706: waveform_sig_rx =-366;
19707: waveform_sig_rx =-384;
19708: waveform_sig_rx =-147;
19709: waveform_sig_rx =-270;
19710: waveform_sig_rx =-322;
19711: waveform_sig_rx =-292;
19712: waveform_sig_rx =-69;
19713: waveform_sig_rx =-375;
19714: waveform_sig_rx =-321;
19715: waveform_sig_rx =-4;
19716: waveform_sig_rx =-331;
19717: waveform_sig_rx =-321;
19718: waveform_sig_rx =-35;
19719: waveform_sig_rx =-204;
19720: waveform_sig_rx =-356;
19721: waveform_sig_rx =-58;
19722: waveform_sig_rx =-120;
19723: waveform_sig_rx =-316;
19724: waveform_sig_rx =-139;
19725: waveform_sig_rx =-52;
19726: waveform_sig_rx =-248;
19727: waveform_sig_rx =-136;
19728: waveform_sig_rx =-171;
19729: waveform_sig_rx =-70;
19730: waveform_sig_rx =-175;
19731: waveform_sig_rx =-89;
19732: waveform_sig_rx =-78;
19733: waveform_sig_rx =-278;
19734: waveform_sig_rx =176;
19735: waveform_sig_rx =-302;
19736: waveform_sig_rx =-71;
19737: waveform_sig_rx =144;
19738: waveform_sig_rx =-328;
19739: waveform_sig_rx =18;
19740: waveform_sig_rx =123;
19741: waveform_sig_rx =-286;
19742: waveform_sig_rx =5;
19743: waveform_sig_rx =137;
19744: waveform_sig_rx =-195;
19745: waveform_sig_rx =6;
19746: waveform_sig_rx =114;
19747: waveform_sig_rx =-35;
19748: waveform_sig_rx =-114;
19749: waveform_sig_rx =150;
19750: waveform_sig_rx =45;
19751: waveform_sig_rx =-56;
19752: waveform_sig_rx =-1;
19753: waveform_sig_rx =237;
19754: waveform_sig_rx =-123;
19755: waveform_sig_rx =0;
19756: waveform_sig_rx =298;
19757: waveform_sig_rx =-91;
19758: waveform_sig_rx =16;
19759: waveform_sig_rx =242;
19760: waveform_sig_rx =35;
19761: waveform_sig_rx =-1;
19762: waveform_sig_rx =171;
19763: waveform_sig_rx =177;
19764: waveform_sig_rx =34;
19765: waveform_sig_rx =83;
19766: waveform_sig_rx =324;
19767: waveform_sig_rx =0;
19768: waveform_sig_rx =143;
19769: waveform_sig_rx =185;
19770: waveform_sig_rx =137;
19771: waveform_sig_rx =156;
19772: waveform_sig_rx =232;
19773: waveform_sig_rx =126;
19774: waveform_sig_rx =115;
19775: waveform_sig_rx =429;
19776: waveform_sig_rx =-67;
19777: waveform_sig_rx =304;
19778: waveform_sig_rx =338;
19779: waveform_sig_rx =-7;
19780: waveform_sig_rx =317;
19781: waveform_sig_rx =387;
19782: waveform_sig_rx =45;
19783: waveform_sig_rx =301;
19784: waveform_sig_rx =410;
19785: waveform_sig_rx =95;
19786: waveform_sig_rx =314;
19787: waveform_sig_rx =360;
19788: waveform_sig_rx =272;
19789: waveform_sig_rx =150;
19790: waveform_sig_rx =435;
19791: waveform_sig_rx =355;
19792: waveform_sig_rx =133;
19793: waveform_sig_rx =364;
19794: waveform_sig_rx =509;
19795: waveform_sig_rx =115;
19796: waveform_sig_rx =419;
19797: waveform_sig_rx =485;
19798: waveform_sig_rx =236;
19799: waveform_sig_rx =333;
19800: waveform_sig_rx =452;
19801: waveform_sig_rx =427;
19802: waveform_sig_rx =244;
19803: waveform_sig_rx =467;
19804: waveform_sig_rx =505;
19805: waveform_sig_rx =222;
19806: waveform_sig_rx =431;
19807: waveform_sig_rx =612;
19808: waveform_sig_rx =231;
19809: waveform_sig_rx =500;
19810: waveform_sig_rx =442;
19811: waveform_sig_rx =424;
19812: waveform_sig_rx =488;
19813: waveform_sig_rx =491;
19814: waveform_sig_rx =398;
19815: waveform_sig_rx =444;
19816: waveform_sig_rx =643;
19817: waveform_sig_rx =263;
19818: waveform_sig_rx =606;
19819: waveform_sig_rx =575;
19820: waveform_sig_rx =322;
19821: waveform_sig_rx =596;
19822: waveform_sig_rx =639;
19823: waveform_sig_rx =345;
19824: waveform_sig_rx =552;
19825: waveform_sig_rx =702;
19826: waveform_sig_rx =382;
19827: waveform_sig_rx =529;
19828: waveform_sig_rx =677;
19829: waveform_sig_rx =549;
19830: waveform_sig_rx =380;
19831: waveform_sig_rx =786;
19832: waveform_sig_rx =579;
19833: waveform_sig_rx =410;
19834: waveform_sig_rx =735;
19835: waveform_sig_rx =687;
19836: waveform_sig_rx =448;
19837: waveform_sig_rx =676;
19838: waveform_sig_rx =684;
19839: waveform_sig_rx =587;
19840: waveform_sig_rx =538;
19841: waveform_sig_rx =762;
19842: waveform_sig_rx =703;
19843: waveform_sig_rx =406;
19844: waveform_sig_rx =824;
19845: waveform_sig_rx =720;
19846: waveform_sig_rx =469;
19847: waveform_sig_rx =763;
19848: waveform_sig_rx =815;
19849: waveform_sig_rx =494;
19850: waveform_sig_rx =783;
19851: waveform_sig_rx =635;
19852: waveform_sig_rx =703;
19853: waveform_sig_rx =752;
19854: waveform_sig_rx =709;
19855: waveform_sig_rx =678;
19856: waveform_sig_rx =713;
19857: waveform_sig_rx =860;
19858: waveform_sig_rx =547;
19859: waveform_sig_rx =831;
19860: waveform_sig_rx =818;
19861: waveform_sig_rx =592;
19862: waveform_sig_rx =795;
19863: waveform_sig_rx =923;
19864: waveform_sig_rx =578;
19865: waveform_sig_rx =766;
19866: waveform_sig_rx =998;
19867: waveform_sig_rx =548;
19868: waveform_sig_rx =800;
19869: waveform_sig_rx =969;
19870: waveform_sig_rx =699;
19871: waveform_sig_rx =699;
19872: waveform_sig_rx =1015;
19873: waveform_sig_rx =749;
19874: waveform_sig_rx =744;
19875: waveform_sig_rx =897;
19876: waveform_sig_rx =925;
19877: waveform_sig_rx =704;
19878: waveform_sig_rx =852;
19879: waveform_sig_rx =962;
19880: waveform_sig_rx =788;
19881: waveform_sig_rx =722;
19882: waveform_sig_rx =1027;
19883: waveform_sig_rx =865;
19884: waveform_sig_rx =659;
19885: waveform_sig_rx =1071;
19886: waveform_sig_rx =893;
19887: waveform_sig_rx =720;
19888: waveform_sig_rx =1004;
19889: waveform_sig_rx =987;
19890: waveform_sig_rx =765;
19891: waveform_sig_rx =1014;
19892: waveform_sig_rx =822;
19893: waveform_sig_rx =977;
19894: waveform_sig_rx =903;
19895: waveform_sig_rx =924;
19896: waveform_sig_rx =903;
19897: waveform_sig_rx =868;
19898: waveform_sig_rx =1080;
19899: waveform_sig_rx =750;
19900: waveform_sig_rx =997;
19901: waveform_sig_rx =1054;
19902: waveform_sig_rx =753;
19903: waveform_sig_rx =997;
19904: waveform_sig_rx =1157;
19905: waveform_sig_rx =702;
19906: waveform_sig_rx =1034;
19907: waveform_sig_rx =1174;
19908: waveform_sig_rx =705;
19909: waveform_sig_rx =1056;
19910: waveform_sig_rx =1113;
19911: waveform_sig_rx =858;
19912: waveform_sig_rx =946;
19913: waveform_sig_rx =1135;
19914: waveform_sig_rx =940;
19915: waveform_sig_rx =939;
19916: waveform_sig_rx =1015;
19917: waveform_sig_rx =1152;
19918: waveform_sig_rx =848;
19919: waveform_sig_rx =1013;
19920: waveform_sig_rx =1199;
19921: waveform_sig_rx =897;
19922: waveform_sig_rx =941;
19923: waveform_sig_rx =1235;
19924: waveform_sig_rx =934;
19925: waveform_sig_rx =891;
19926: waveform_sig_rx =1198;
19927: waveform_sig_rx =997;
19928: waveform_sig_rx =919;
19929: waveform_sig_rx =1109;
19930: waveform_sig_rx =1114;
19931: waveform_sig_rx =921;
19932: waveform_sig_rx =1110;
19933: waveform_sig_rx =973;
19934: waveform_sig_rx =1124;
19935: waveform_sig_rx =999;
19936: waveform_sig_rx =1111;
19937: waveform_sig_rx =1012;
19938: waveform_sig_rx =995;
19939: waveform_sig_rx =1275;
19940: waveform_sig_rx =838;
19941: waveform_sig_rx =1153;
19942: waveform_sig_rx =1227;
19943: waveform_sig_rx =817;
19944: waveform_sig_rx =1235;
19945: waveform_sig_rx =1246;
19946: waveform_sig_rx =783;
19947: waveform_sig_rx =1259;
19948: waveform_sig_rx =1214;
19949: waveform_sig_rx =860;
19950: waveform_sig_rx =1219;
19951: waveform_sig_rx =1154;
19952: waveform_sig_rx =1013;
19953: waveform_sig_rx =1016;
19954: waveform_sig_rx =1209;
19955: waveform_sig_rx =1087;
19956: waveform_sig_rx =999;
19957: waveform_sig_rx =1146;
19958: waveform_sig_rx =1264;
19959: waveform_sig_rx =904;
19960: waveform_sig_rx =1200;
19961: waveform_sig_rx =1267;
19962: waveform_sig_rx =969;
19963: waveform_sig_rx =1102;
19964: waveform_sig_rx =1297;
19965: waveform_sig_rx =1059;
19966: waveform_sig_rx =1022;
19967: waveform_sig_rx =1291;
19968: waveform_sig_rx =1145;
19969: waveform_sig_rx =1032;
19970: waveform_sig_rx =1204;
19971: waveform_sig_rx =1257;
19972: waveform_sig_rx =1009;
19973: waveform_sig_rx =1207;
19974: waveform_sig_rx =1093;
19975: waveform_sig_rx =1208;
19976: waveform_sig_rx =1074;
19977: waveform_sig_rx =1250;
19978: waveform_sig_rx =1036;
19979: waveform_sig_rx =1111;
19980: waveform_sig_rx =1340;
19981: waveform_sig_rx =865;
19982: waveform_sig_rx =1312;
19983: waveform_sig_rx =1224;
19984: waveform_sig_rx =890;
19985: waveform_sig_rx =1366;
19986: waveform_sig_rx =1193;
19987: waveform_sig_rx =935;
19988: waveform_sig_rx =1311;
19989: waveform_sig_rx =1204;
19990: waveform_sig_rx =1009;
19991: waveform_sig_rx =1203;
19992: waveform_sig_rx =1239;
19993: waveform_sig_rx =1096;
19994: waveform_sig_rx =1007;
19995: waveform_sig_rx =1331;
19996: waveform_sig_rx =1094;
19997: waveform_sig_rx =1016;
19998: waveform_sig_rx =1243;
19999: waveform_sig_rx =1239;
20000: waveform_sig_rx =956;
20001: waveform_sig_rx =1232;
20002: waveform_sig_rx =1280;
20003: waveform_sig_rx =1003;
20004: waveform_sig_rx =1158;
20005: waveform_sig_rx =1298;
20006: waveform_sig_rx =1074;
20007: waveform_sig_rx =1067;
20008: waveform_sig_rx =1254;
20009: waveform_sig_rx =1164;
20010: waveform_sig_rx =1009;
20011: waveform_sig_rx =1190;
20012: waveform_sig_rx =1318;
20013: waveform_sig_rx =925;
20014: waveform_sig_rx =1242;
20015: waveform_sig_rx =1116;
20016: waveform_sig_rx =1133;
20017: waveform_sig_rx =1141;
20018: waveform_sig_rx =1243;
20019: waveform_sig_rx =1002;
20020: waveform_sig_rx =1223;
20021: waveform_sig_rx =1264;
20022: waveform_sig_rx =884;
20023: waveform_sig_rx =1364;
20024: waveform_sig_rx =1125;
20025: waveform_sig_rx =979;
20026: waveform_sig_rx =1295;
20027: waveform_sig_rx =1174;
20028: waveform_sig_rx =953;
20029: waveform_sig_rx =1239;
20030: waveform_sig_rx =1227;
20031: waveform_sig_rx =972;
20032: waveform_sig_rx =1174;
20033: waveform_sig_rx =1271;
20034: waveform_sig_rx =1024;
20035: waveform_sig_rx =1039;
20036: waveform_sig_rx =1327;
20037: waveform_sig_rx =1047;
20038: waveform_sig_rx =1015;
20039: waveform_sig_rx =1214;
20040: waveform_sig_rx =1214;
20041: waveform_sig_rx =908;
20042: waveform_sig_rx =1248;
20043: waveform_sig_rx =1179;
20044: waveform_sig_rx =970;
20045: waveform_sig_rx =1118;
20046: waveform_sig_rx =1203;
20047: waveform_sig_rx =1094;
20048: waveform_sig_rx =967;
20049: waveform_sig_rx =1232;
20050: waveform_sig_rx =1158;
20051: waveform_sig_rx =871;
20052: waveform_sig_rx =1261;
20053: waveform_sig_rx =1172;
20054: waveform_sig_rx =870;
20055: waveform_sig_rx =1278;
20056: waveform_sig_rx =923;
20057: waveform_sig_rx =1162;
20058: waveform_sig_rx =1054;
20059: waveform_sig_rx =1079;
20060: waveform_sig_rx =998;
20061: waveform_sig_rx =1094;
20062: waveform_sig_rx =1146;
20063: waveform_sig_rx =858;
20064: waveform_sig_rx =1187;
20065: waveform_sig_rx =1069;
20066: waveform_sig_rx =860;
20067: waveform_sig_rx =1193;
20068: waveform_sig_rx =1086;
20069: waveform_sig_rx =826;
20070: waveform_sig_rx =1128;
20071: waveform_sig_rx =1104;
20072: waveform_sig_rx =865;
20073: waveform_sig_rx =1058;
20074: waveform_sig_rx =1170;
20075: waveform_sig_rx =878;
20076: waveform_sig_rx =936;
20077: waveform_sig_rx =1236;
20078: waveform_sig_rx =865;
20079: waveform_sig_rx =957;
20080: waveform_sig_rx =1097;
20081: waveform_sig_rx =1037;
20082: waveform_sig_rx =869;
20083: waveform_sig_rx =1075;
20084: waveform_sig_rx =1078;
20085: waveform_sig_rx =880;
20086: waveform_sig_rx =943;
20087: waveform_sig_rx =1139;
20088: waveform_sig_rx =930;
20089: waveform_sig_rx =831;
20090: waveform_sig_rx =1204;
20091: waveform_sig_rx =928;
20092: waveform_sig_rx =772;
20093: waveform_sig_rx =1151;
20094: waveform_sig_rx =943;
20095: waveform_sig_rx =812;
20096: waveform_sig_rx =1096;
20097: waveform_sig_rx =769;
20098: waveform_sig_rx =1079;
20099: waveform_sig_rx =841;
20100: waveform_sig_rx =983;
20101: waveform_sig_rx =833;
20102: waveform_sig_rx =908;
20103: waveform_sig_rx =1013;
20104: waveform_sig_rx =678;
20105: waveform_sig_rx =1058;
20106: waveform_sig_rx =922;
20107: waveform_sig_rx =701;
20108: waveform_sig_rx =1050;
20109: waveform_sig_rx =915;
20110: waveform_sig_rx =674;
20111: waveform_sig_rx =990;
20112: waveform_sig_rx =974;
20113: waveform_sig_rx =651;
20114: waveform_sig_rx =911;
20115: waveform_sig_rx =1003;
20116: waveform_sig_rx =620;
20117: waveform_sig_rx =859;
20118: waveform_sig_rx =988;
20119: waveform_sig_rx =692;
20120: waveform_sig_rx =829;
20121: waveform_sig_rx =820;
20122: waveform_sig_rx =919;
20123: waveform_sig_rx =643;
20124: waveform_sig_rx =858;
20125: waveform_sig_rx =950;
20126: waveform_sig_rx =612;
20127: waveform_sig_rx =822;
20128: waveform_sig_rx =978;
20129: waveform_sig_rx =663;
20130: waveform_sig_rx =725;
20131: waveform_sig_rx =947;
20132: waveform_sig_rx =728;
20133: waveform_sig_rx =638;
20134: waveform_sig_rx =914;
20135: waveform_sig_rx =774;
20136: waveform_sig_rx =628;
20137: waveform_sig_rx =864;
20138: waveform_sig_rx =603;
20139: waveform_sig_rx =859;
20140: waveform_sig_rx =625;
20141: waveform_sig_rx =828;
20142: waveform_sig_rx =609;
20143: waveform_sig_rx =733;
20144: waveform_sig_rx =834;
20145: waveform_sig_rx =468;
20146: waveform_sig_rx =854;
20147: waveform_sig_rx =723;
20148: waveform_sig_rx =451;
20149: waveform_sig_rx =892;
20150: waveform_sig_rx =701;
20151: waveform_sig_rx =405;
20152: waveform_sig_rx =862;
20153: waveform_sig_rx =671;
20154: waveform_sig_rx =453;
20155: waveform_sig_rx =787;
20156: waveform_sig_rx =689;
20157: waveform_sig_rx =476;
20158: waveform_sig_rx =623;
20159: waveform_sig_rx =713;
20160: waveform_sig_rx =539;
20161: waveform_sig_rx =540;
20162: waveform_sig_rx =638;
20163: waveform_sig_rx =699;
20164: waveform_sig_rx =347;
20165: waveform_sig_rx =696;
20166: waveform_sig_rx =673;
20167: waveform_sig_rx =363;
20168: waveform_sig_rx =615;
20169: waveform_sig_rx =695;
20170: waveform_sig_rx =409;
20171: waveform_sig_rx =482;
20172: waveform_sig_rx =680;
20173: waveform_sig_rx =460;
20174: waveform_sig_rx =414;
20175: waveform_sig_rx =625;
20176: waveform_sig_rx =528;
20177: waveform_sig_rx =388;
20178: waveform_sig_rx =560;
20179: waveform_sig_rx =386;
20180: waveform_sig_rx =573;
20181: waveform_sig_rx =365;
20182: waveform_sig_rx =604;
20183: waveform_sig_rx =293;
20184: waveform_sig_rx =523;
20185: waveform_sig_rx =544;
20186: waveform_sig_rx =170;
20187: waveform_sig_rx =638;
20188: waveform_sig_rx =391;
20189: waveform_sig_rx =179;
20190: waveform_sig_rx =661;
20191: waveform_sig_rx =361;
20192: waveform_sig_rx =197;
20193: waveform_sig_rx =590;
20194: waveform_sig_rx =349;
20195: waveform_sig_rx =219;
20196: waveform_sig_rx =465;
20197: waveform_sig_rx =404;
20198: waveform_sig_rx =230;
20199: waveform_sig_rx =294;
20200: waveform_sig_rx =464;
20201: waveform_sig_rx =258;
20202: waveform_sig_rx =235;
20203: waveform_sig_rx =440;
20204: waveform_sig_rx =387;
20205: waveform_sig_rx =88;
20206: waveform_sig_rx =463;
20207: waveform_sig_rx =347;
20208: waveform_sig_rx =102;
20209: waveform_sig_rx =363;
20210: waveform_sig_rx =373;
20211: waveform_sig_rx =159;
20212: waveform_sig_rx =225;
20213: waveform_sig_rx =363;
20214: waveform_sig_rx =195;
20215: waveform_sig_rx =88;
20216: waveform_sig_rx =338;
20217: waveform_sig_rx =267;
20218: waveform_sig_rx =33;
20219: waveform_sig_rx =306;
20220: waveform_sig_rx =111;
20221: waveform_sig_rx =228;
20222: waveform_sig_rx =121;
20223: waveform_sig_rx =267;
20224: waveform_sig_rx =-37;
20225: waveform_sig_rx =298;
20226: waveform_sig_rx =172;
20227: waveform_sig_rx =-77;
20228: waveform_sig_rx =358;
20229: waveform_sig_rx =39;
20230: waveform_sig_rx =-21;
20231: waveform_sig_rx =318;
20232: waveform_sig_rx =77;
20233: waveform_sig_rx =-60;
20234: waveform_sig_rx =263;
20235: waveform_sig_rx =79;
20236: waveform_sig_rx =-52;
20237: waveform_sig_rx =153;
20238: waveform_sig_rx =122;
20239: waveform_sig_rx =-66;
20240: waveform_sig_rx =5;
20241: waveform_sig_rx =208;
20242: waveform_sig_rx =-73;
20243: waveform_sig_rx =-94;
20244: waveform_sig_rx =187;
20245: waveform_sig_rx =1;
20246: waveform_sig_rx =-181;
20247: waveform_sig_rx =177;
20248: waveform_sig_rx =-29;
20249: waveform_sig_rx =-130;
20250: waveform_sig_rx =1;
20251: waveform_sig_rx =63;
20252: waveform_sig_rx =-117;
20253: waveform_sig_rx =-160;
20254: waveform_sig_rx =123;
20255: waveform_sig_rx =-115;
20256: waveform_sig_rx =-238;
20257: waveform_sig_rx =109;
20258: waveform_sig_rx =-95;
20259: waveform_sig_rx =-239;
20260: waveform_sig_rx =33;
20261: waveform_sig_rx =-236;
20262: waveform_sig_rx =-24;
20263: waveform_sig_rx =-170;
20264: waveform_sig_rx =-67;
20265: waveform_sig_rx =-302;
20266: waveform_sig_rx =16;
20267: waveform_sig_rx =-173;
20268: waveform_sig_rx =-335;
20269: waveform_sig_rx =37;
20270: waveform_sig_rx =-259;
20271: waveform_sig_rx =-288;
20272: waveform_sig_rx =-22;
20273: waveform_sig_rx =-215;
20274: waveform_sig_rx =-371;
20275: waveform_sig_rx =-76;
20276: waveform_sig_rx =-208;
20277: waveform_sig_rx =-417;
20278: waveform_sig_rx =-146;
20279: waveform_sig_rx =-130;
20280: waveform_sig_rx =-454;
20281: waveform_sig_rx =-250;
20282: waveform_sig_rx =-98;
20283: waveform_sig_rx =-433;
20284: waveform_sig_rx =-335;
20285: waveform_sig_rx =-172;
20286: waveform_sig_rx =-333;
20287: waveform_sig_rx =-447;
20288: waveform_sig_rx =-203;
20289: waveform_sig_rx =-300;
20290: waveform_sig_rx =-437;
20291: waveform_sig_rx =-347;
20292: waveform_sig_rx =-184;
20293: waveform_sig_rx =-483;
20294: waveform_sig_rx =-439;
20295: waveform_sig_rx =-140;
20296: waveform_sig_rx =-479;
20297: waveform_sig_rx =-495;
20298: waveform_sig_rx =-185;
20299: waveform_sig_rx =-432;
20300: waveform_sig_rx =-491;
20301: waveform_sig_rx =-276;
20302: waveform_sig_rx =-533;
20303: waveform_sig_rx =-289;
20304: waveform_sig_rx =-483;
20305: waveform_sig_rx =-376;
20306: waveform_sig_rx =-574;
20307: waveform_sig_rx =-336;
20308: waveform_sig_rx =-479;
20309: waveform_sig_rx =-602;
20310: waveform_sig_rx =-322;
20311: waveform_sig_rx =-512;
20312: waveform_sig_rx =-620;
20313: waveform_sig_rx =-321;
20314: waveform_sig_rx =-488;
20315: waveform_sig_rx =-732;
20316: waveform_sig_rx =-299;
20317: waveform_sig_rx =-524;
20318: waveform_sig_rx =-737;
20319: waveform_sig_rx =-378;
20320: waveform_sig_rx =-496;
20321: waveform_sig_rx =-745;
20322: waveform_sig_rx =-483;
20323: waveform_sig_rx =-445;
20324: waveform_sig_rx =-689;
20325: waveform_sig_rx =-606;
20326: waveform_sig_rx =-491;
20327: waveform_sig_rx =-588;
20328: waveform_sig_rx =-733;
20329: waveform_sig_rx =-496;
20330: waveform_sig_rx =-538;
20331: waveform_sig_rx =-748;
20332: waveform_sig_rx =-618;
20333: waveform_sig_rx =-434;
20334: waveform_sig_rx =-836;
20335: waveform_sig_rx =-664;
20336: waveform_sig_rx =-444;
20337: waveform_sig_rx =-830;
20338: waveform_sig_rx =-696;
20339: waveform_sig_rx =-515;
20340: waveform_sig_rx =-731;
20341: waveform_sig_rx =-729;
20342: waveform_sig_rx =-630;
20343: waveform_sig_rx =-782;
20344: waveform_sig_rx =-577;
20345: waveform_sig_rx =-821;
20346: waveform_sig_rx =-611;
20347: waveform_sig_rx =-847;
20348: waveform_sig_rx =-616;
20349: waveform_sig_rx =-707;
20350: waveform_sig_rx =-907;
20351: waveform_sig_rx =-547;
20352: waveform_sig_rx =-756;
20353: waveform_sig_rx =-961;
20354: waveform_sig_rx =-521;
20355: waveform_sig_rx =-783;
20356: waveform_sig_rx =-1026;
20357: waveform_sig_rx =-495;
20358: waveform_sig_rx =-856;
20359: waveform_sig_rx =-952;
20360: waveform_sig_rx =-606;
20361: waveform_sig_rx =-800;
20362: waveform_sig_rx =-942;
20363: waveform_sig_rx =-763;
20364: waveform_sig_rx =-716;
20365: waveform_sig_rx =-917;
20366: waveform_sig_rx =-907;
20367: waveform_sig_rx =-715;
20368: waveform_sig_rx =-823;
20369: waveform_sig_rx =-998;
20370: waveform_sig_rx =-687;
20371: waveform_sig_rx =-780;
20372: waveform_sig_rx =-1042;
20373: waveform_sig_rx =-785;
20374: waveform_sig_rx =-693;
20375: waveform_sig_rx =-1085;
20376: waveform_sig_rx =-810;
20377: waveform_sig_rx =-730;
20378: waveform_sig_rx =-1009;
20379: waveform_sig_rx =-886;
20380: waveform_sig_rx =-793;
20381: waveform_sig_rx =-886;
20382: waveform_sig_rx =-972;
20383: waveform_sig_rx =-873;
20384: waveform_sig_rx =-944;
20385: waveform_sig_rx =-856;
20386: waveform_sig_rx =-991;
20387: waveform_sig_rx =-806;
20388: waveform_sig_rx =-1130;
20389: waveform_sig_rx =-770;
20390: waveform_sig_rx =-951;
20391: waveform_sig_rx =-1144;
20392: waveform_sig_rx =-716;
20393: waveform_sig_rx =-1059;
20394: waveform_sig_rx =-1131;
20395: waveform_sig_rx =-685;
20396: waveform_sig_rx =-1065;
20397: waveform_sig_rx =-1148;
20398: waveform_sig_rx =-663;
20399: waveform_sig_rx =-1124;
20400: waveform_sig_rx =-1086;
20401: waveform_sig_rx =-829;
20402: waveform_sig_rx =-1029;
20403: waveform_sig_rx =-1088;
20404: waveform_sig_rx =-982;
20405: waveform_sig_rx =-891;
20406: waveform_sig_rx =-1088;
20407: waveform_sig_rx =-1122;
20408: waveform_sig_rx =-836;
20409: waveform_sig_rx =-1054;
20410: waveform_sig_rx =-1201;
20411: waveform_sig_rx =-835;
20412: waveform_sig_rx =-1053;
20413: waveform_sig_rx =-1197;
20414: waveform_sig_rx =-932;
20415: waveform_sig_rx =-937;
20416: waveform_sig_rx =-1194;
20417: waveform_sig_rx =-1019;
20418: waveform_sig_rx =-911;
20419: waveform_sig_rx =-1145;
20420: waveform_sig_rx =-1127;
20421: waveform_sig_rx =-938;
20422: waveform_sig_rx =-1058;
20423: waveform_sig_rx =-1157;
20424: waveform_sig_rx =-1007;
20425: waveform_sig_rx =-1110;
20426: waveform_sig_rx =-1037;
20427: waveform_sig_rx =-1104;
20428: waveform_sig_rx =-973;
20429: waveform_sig_rx =-1295;
20430: waveform_sig_rx =-866;
20431: waveform_sig_rx =-1166;
20432: waveform_sig_rx =-1229;
20433: waveform_sig_rx =-824;
20434: waveform_sig_rx =-1275;
20435: waveform_sig_rx =-1178;
20436: waveform_sig_rx =-860;
20437: waveform_sig_rx =-1263;
20438: waveform_sig_rx =-1202;
20439: waveform_sig_rx =-913;
20440: waveform_sig_rx =-1220;
20441: waveform_sig_rx =-1190;
20442: waveform_sig_rx =-1044;
20443: waveform_sig_rx =-1066;
20444: waveform_sig_rx =-1281;
20445: waveform_sig_rx =-1110;
20446: waveform_sig_rx =-970;
20447: waveform_sig_rx =-1265;
20448: waveform_sig_rx =-1181;
20449: waveform_sig_rx =-943;
20450: waveform_sig_rx =-1206;
20451: waveform_sig_rx =-1261;
20452: waveform_sig_rx =-958;
20453: waveform_sig_rx =-1187;
20454: waveform_sig_rx =-1245;
20455: waveform_sig_rx =-1053;
20456: waveform_sig_rx =-1064;
20457: waveform_sig_rx =-1276;
20458: waveform_sig_rx =-1149;
20459: waveform_sig_rx =-1020;
20460: waveform_sig_rx =-1238;
20461: waveform_sig_rx =-1260;
20462: waveform_sig_rx =-968;
20463: waveform_sig_rx =-1197;
20464: waveform_sig_rx =-1262;
20465: waveform_sig_rx =-1027;
20466: waveform_sig_rx =-1252;
20467: waveform_sig_rx =-1109;
20468: waveform_sig_rx =-1153;
20469: waveform_sig_rx =-1117;
20470: waveform_sig_rx =-1326;
20471: waveform_sig_rx =-930;
20472: waveform_sig_rx =-1314;
20473: waveform_sig_rx =-1203;
20474: waveform_sig_rx =-961;
20475: waveform_sig_rx =-1331;
20476: waveform_sig_rx =-1168;
20477: waveform_sig_rx =-1005;
20478: waveform_sig_rx =-1260;
20479: waveform_sig_rx =-1270;
20480: waveform_sig_rx =-996;
20481: waveform_sig_rx =-1217;
20482: waveform_sig_rx =-1269;
20483: waveform_sig_rx =-1028;
20484: waveform_sig_rx =-1084;
20485: waveform_sig_rx =-1364;
20486: waveform_sig_rx =-1067;
20487: waveform_sig_rx =-1045;
20488: waveform_sig_rx =-1307;
20489: waveform_sig_rx =-1173;
20490: waveform_sig_rx =-1009;
20491: waveform_sig_rx =-1214;
20492: waveform_sig_rx =-1250;
20493: waveform_sig_rx =-975;
20494: waveform_sig_rx =-1207;
20495: waveform_sig_rx =-1244;
20496: waveform_sig_rx =-1084;
20497: waveform_sig_rx =-1062;
20498: waveform_sig_rx =-1254;
20499: waveform_sig_rx =-1184;
20500: waveform_sig_rx =-953;
20501: waveform_sig_rx =-1276;
20502: waveform_sig_rx =-1261;
20503: waveform_sig_rx =-903;
20504: waveform_sig_rx =-1300;
20505: waveform_sig_rx =-1178;
20506: waveform_sig_rx =-1041;
20507: waveform_sig_rx =-1301;
20508: waveform_sig_rx =-1006;
20509: waveform_sig_rx =-1208;
20510: waveform_sig_rx =-1090;
20511: waveform_sig_rx =-1258;
20512: waveform_sig_rx =-983;
20513: waveform_sig_rx =-1234;
20514: waveform_sig_rx =-1214;
20515: waveform_sig_rx =-955;
20516: waveform_sig_rx =-1241;
20517: waveform_sig_rx =-1218;
20518: waveform_sig_rx =-913;
20519: waveform_sig_rx =-1260;
20520: waveform_sig_rx =-1237;
20521: waveform_sig_rx =-915;
20522: waveform_sig_rx =-1223;
20523: waveform_sig_rx =-1220;
20524: waveform_sig_rx =-1006;
20525: waveform_sig_rx =-1066;
20526: waveform_sig_rx =-1332;
20527: waveform_sig_rx =-993;
20528: waveform_sig_rx =-1030;
20529: waveform_sig_rx =-1275;
20530: waveform_sig_rx =-1077;
20531: waveform_sig_rx =-1001;
20532: waveform_sig_rx =-1174;
20533: waveform_sig_rx =-1154;
20534: waveform_sig_rx =-983;
20535: waveform_sig_rx =-1084;
20536: waveform_sig_rx =-1229;
20537: waveform_sig_rx =-1004;
20538: waveform_sig_rx =-952;
20539: waveform_sig_rx =-1300;
20540: waveform_sig_rx =-1032;
20541: waveform_sig_rx =-888;
20542: waveform_sig_rx =-1260;
20543: waveform_sig_rx =-1063;
20544: waveform_sig_rx =-885;
20545: waveform_sig_rx =-1193;
20546: waveform_sig_rx =-1017;
20547: waveform_sig_rx =-1064;
20548: waveform_sig_rx =-1098;
20549: waveform_sig_rx =-947;
20550: waveform_sig_rx =-1141;
20551: waveform_sig_rx =-947;
20552: waveform_sig_rx =-1211;
20553: waveform_sig_rx =-852;
20554: waveform_sig_rx =-1136;
20555: waveform_sig_rx =-1134;
20556: waveform_sig_rx =-822;
20557: waveform_sig_rx =-1183;
20558: waveform_sig_rx =-1094;
20559: waveform_sig_rx =-798;
20560: waveform_sig_rx =-1149;
20561: waveform_sig_rx =-1116;
20562: waveform_sig_rx =-776;
20563: waveform_sig_rx =-1126;
20564: waveform_sig_rx =-1108;
20565: waveform_sig_rx =-842;
20566: waveform_sig_rx =-1003;
20567: waveform_sig_rx =-1210;
20568: waveform_sig_rx =-793;
20569: waveform_sig_rx =-987;
20570: waveform_sig_rx =-1060;
20571: waveform_sig_rx =-959;
20572: waveform_sig_rx =-881;
20573: waveform_sig_rx =-964;
20574: waveform_sig_rx =-1116;
20575: waveform_sig_rx =-774;
20576: waveform_sig_rx =-946;
20577: waveform_sig_rx =-1148;
20578: waveform_sig_rx =-758;
20579: waveform_sig_rx =-885;
20580: waveform_sig_rx =-1130;
20581: waveform_sig_rx =-828;
20582: waveform_sig_rx =-834;
20583: waveform_sig_rx =-1024;
20584: waveform_sig_rx =-935;
20585: waveform_sig_rx =-738;
20586: waveform_sig_rx =-981;
20587: waveform_sig_rx =-886;
20588: waveform_sig_rx =-882;
20589: waveform_sig_rx =-923;
20590: waveform_sig_rx =-818;
20591: waveform_sig_rx =-935;
20592: waveform_sig_rx =-766;
20593: waveform_sig_rx =-1065;
20594: waveform_sig_rx =-669;
20595: waveform_sig_rx =-985;
20596: waveform_sig_rx =-953;
20597: waveform_sig_rx =-614;
20598: waveform_sig_rx =-1019;
20599: waveform_sig_rx =-899;
20600: waveform_sig_rx =-579;
20601: waveform_sig_rx =-1026;
20602: waveform_sig_rx =-904;
20603: waveform_sig_rx =-580;
20604: waveform_sig_rx =-1012;
20605: waveform_sig_rx =-848;
20606: waveform_sig_rx =-654;
20607: waveform_sig_rx =-838;
20608: waveform_sig_rx =-924;
20609: waveform_sig_rx =-679;
20610: waveform_sig_rx =-768;
20611: waveform_sig_rx =-836;
20612: waveform_sig_rx =-847;
20613: waveform_sig_rx =-587;
20614: waveform_sig_rx =-843;
20615: waveform_sig_rx =-912;
20616: waveform_sig_rx =-504;
20617: waveform_sig_rx =-864;
20618: waveform_sig_rx =-853;
20619: waveform_sig_rx =-578;
20620: waveform_sig_rx =-725;
20621: waveform_sig_rx =-854;
20622: waveform_sig_rx =-667;
20623: waveform_sig_rx =-614;
20624: waveform_sig_rx =-835;
20625: waveform_sig_rx =-731;
20626: waveform_sig_rx =-526;
20627: waveform_sig_rx =-801;
20628: waveform_sig_rx =-665;
20629: waveform_sig_rx =-674;
20630: waveform_sig_rx =-670;
20631: waveform_sig_rx =-626;
20632: waveform_sig_rx =-679;
20633: waveform_sig_rx =-562;
20634: waveform_sig_rx =-846;
20635: waveform_sig_rx =-365;
20636: waveform_sig_rx =-795;
20637: waveform_sig_rx =-707;
20638: waveform_sig_rx =-360;
20639: waveform_sig_rx =-874;
20640: waveform_sig_rx =-581;
20641: waveform_sig_rx =-375;
20642: waveform_sig_rx =-827;
20643: waveform_sig_rx =-562;
20644: waveform_sig_rx =-412;
20645: waveform_sig_rx =-721;
20646: waveform_sig_rx =-590;
20647: waveform_sig_rx =-473;
20648: waveform_sig_rx =-549;
20649: waveform_sig_rx =-714;
20650: waveform_sig_rx =-438;
20651: waveform_sig_rx =-483;
20652: waveform_sig_rx =-656;
20653: waveform_sig_rx =-560;
20654: waveform_sig_rx =-333;
20655: waveform_sig_rx =-649;
20656: waveform_sig_rx =-575;
20657: waveform_sig_rx =-277;
20658: waveform_sig_rx =-604;
20659: waveform_sig_rx =-548;
20660: waveform_sig_rx =-345;
20661: waveform_sig_rx =-474;
20662: waveform_sig_rx =-571;
20663: waveform_sig_rx =-436;
20664: waveform_sig_rx =-363;
20665: waveform_sig_rx =-578;
20666: waveform_sig_rx =-497;
20667: waveform_sig_rx =-244;
20668: waveform_sig_rx =-565;
20669: waveform_sig_rx =-439;
20670: waveform_sig_rx =-388;
20671: waveform_sig_rx =-458;
20672: waveform_sig_rx =-387;
20673: waveform_sig_rx =-397;
20674: waveform_sig_rx =-380;
20675: waveform_sig_rx =-556;
20676: waveform_sig_rx =-119;
20677: waveform_sig_rx =-597;
20678: waveform_sig_rx =-341;
20679: waveform_sig_rx =-169;
20680: waveform_sig_rx =-615;
20681: waveform_sig_rx =-256;
20682: waveform_sig_rx =-201;
20683: waveform_sig_rx =-523;
20684: waveform_sig_rx =-310;
20685: waveform_sig_rx =-185;
20686: waveform_sig_rx =-414;
20687: waveform_sig_rx =-349;
20688: waveform_sig_rx =-186;
20689: waveform_sig_rx =-267;
20690: waveform_sig_rx =-485;
20691: waveform_sig_rx =-123;
20692: waveform_sig_rx =-228;
20693: waveform_sig_rx =-404;
20694: waveform_sig_rx =-235;
20695: waveform_sig_rx =-104;
20696: waveform_sig_rx =-391;
20697: waveform_sig_rx =-261;
20698: waveform_sig_rx =-69;
20699: waveform_sig_rx =-303;
20700: waveform_sig_rx =-261;
20701: waveform_sig_rx =-106;
20702: waveform_sig_rx =-151;
20703: waveform_sig_rx =-337;
20704: waveform_sig_rx =-134;
20705: waveform_sig_rx =-29;
20706: waveform_sig_rx =-346;
20707: waveform_sig_rx =-179;
20708: waveform_sig_rx =51;
20709: waveform_sig_rx =-317;
20710: waveform_sig_rx =-106;
20711: waveform_sig_rx =-129;
20712: waveform_sig_rx =-189;
20713: waveform_sig_rx =-72;
20714: waveform_sig_rx =-117;
20715: waveform_sig_rx =-118;
20716: waveform_sig_rx =-196;
20717: waveform_sig_rx =120;
20718: waveform_sig_rx =-299;
20719: waveform_sig_rx =-30;
20720: waveform_sig_rx =55;
20721: waveform_sig_rx =-248;
20722: waveform_sig_rx =-16;
20723: waveform_sig_rx =93;
20724: waveform_sig_rx =-176;
20725: waveform_sig_rx =-92;
20726: waveform_sig_rx =170;
20727: waveform_sig_rx =-148;
20728: waveform_sig_rx =-68;
20729: waveform_sig_rx =155;
20730: waveform_sig_rx =-15;
20731: waveform_sig_rx =-207;
20732: waveform_sig_rx =217;
20733: waveform_sig_rx =22;
20734: waveform_sig_rx =-108;
20735: waveform_sig_rx =80;
20736: waveform_sig_rx =137;
20737: waveform_sig_rx =-57;
20738: waveform_sig_rx =31;
20739: waveform_sig_rx =199;
20740: waveform_sig_rx =35;
20741: waveform_sig_rx =-38;
20742: waveform_sig_rx =212;
20743: waveform_sig_rx =170;
20744: waveform_sig_rx =-104;
20745: waveform_sig_rx =209;
20746: waveform_sig_rx =228;
20747: waveform_sig_rx =-65;
20748: waveform_sig_rx =173;
20749: waveform_sig_rx =310;
20750: waveform_sig_rx =-36;
20751: waveform_sig_rx =222;
20752: waveform_sig_rx =124;
20753: waveform_sig_rx =120;
20754: waveform_sig_rx =232;
20755: waveform_sig_rx =140;
20756: waveform_sig_rx =209;
20757: waveform_sig_rx =114;
20758: waveform_sig_rx =366;
20759: waveform_sig_rx =43;
20760: waveform_sig_rx =234;
20761: waveform_sig_rx =340;
20762: waveform_sig_rx =83;
20763: waveform_sig_rx =220;
20764: waveform_sig_rx =448;
20765: waveform_sig_rx =70;
20766: waveform_sig_rx =184;
20767: waveform_sig_rx =511;
20768: waveform_sig_rx =57;
20769: waveform_sig_rx =267;
20770: waveform_sig_rx =438;
20771: waveform_sig_rx =209;
20772: waveform_sig_rx =159;
20773: waveform_sig_rx =447;
20774: waveform_sig_rx =299;
20775: waveform_sig_rx =222;
20776: waveform_sig_rx =351;
20777: waveform_sig_rx =458;
20778: waveform_sig_rx =224;
20779: waveform_sig_rx =325;
20780: waveform_sig_rx =477;
20781: waveform_sig_rx =314;
20782: waveform_sig_rx =250;
20783: waveform_sig_rx =506;
20784: waveform_sig_rx =440;
20785: waveform_sig_rx =157;
20786: waveform_sig_rx =562;
20787: waveform_sig_rx =471;
20788: waveform_sig_rx =224;
20789: waveform_sig_rx =517;
20790: waveform_sig_rx =509;
20791: waveform_sig_rx =312;
20792: waveform_sig_rx =499;
20793: waveform_sig_rx =372;
20794: waveform_sig_rx =490;
20795: waveform_sig_rx =450;
20796: waveform_sig_rx =441;
20797: waveform_sig_rx =505;
20798: waveform_sig_rx =333;
20799: waveform_sig_rx =674;
20800: waveform_sig_rx =316;
20801: waveform_sig_rx =480;
20802: waveform_sig_rx =691;
20803: waveform_sig_rx =298;
20804: waveform_sig_rx =540;
20805: waveform_sig_rx =744;
20806: waveform_sig_rx =271;
20807: waveform_sig_rx =539;
20808: waveform_sig_rx =729;
20809: waveform_sig_rx =318;
20810: waveform_sig_rx =565;
20811: waveform_sig_rx =659;
20812: waveform_sig_rx =485;
20813: waveform_sig_rx =449;
20814: waveform_sig_rx =721;
20815: waveform_sig_rx =587;
20816: waveform_sig_rx =484;
20817: waveform_sig_rx =615;
20818: waveform_sig_rx =750;
20819: waveform_sig_rx =436;
20820: waveform_sig_rx =586;
20821: waveform_sig_rx =796;
20822: waveform_sig_rx =528;
20823: waveform_sig_rx =527;
20824: waveform_sig_rx =858;
20825: waveform_sig_rx =626;
20826: waveform_sig_rx =500;
20827: waveform_sig_rx =841;
20828: waveform_sig_rx =676;
20829: waveform_sig_rx =569;
20830: waveform_sig_rx =714;
20831: waveform_sig_rx =773;
20832: waveform_sig_rx =601;
20833: waveform_sig_rx =674;
20834: waveform_sig_rx =668;
20835: waveform_sig_rx =736;
20836: waveform_sig_rx =641;
20837: waveform_sig_rx =780;
20838: waveform_sig_rx =673;
20839: waveform_sig_rx =615;
20840: waveform_sig_rx =975;
20841: waveform_sig_rx =477;
20842: waveform_sig_rx =793;
20843: waveform_sig_rx =888;
20844: waveform_sig_rx =490;
20845: waveform_sig_rx =856;
20846: waveform_sig_rx =908;
20847: waveform_sig_rx =516;
20848: waveform_sig_rx =820;
20849: waveform_sig_rx =947;
20850: waveform_sig_rx =573;
20851: waveform_sig_rx =858;
20852: waveform_sig_rx =883;
20853: waveform_sig_rx =745;
20854: waveform_sig_rx =689;
20855: waveform_sig_rx =930;
20856: waveform_sig_rx =826;
20857: waveform_sig_rx =691;
20858: waveform_sig_rx =841;
20859: waveform_sig_rx =1010;
20860: waveform_sig_rx =606;
20861: waveform_sig_rx =864;
20862: waveform_sig_rx =1020;
20863: waveform_sig_rx =682;
20864: waveform_sig_rx =849;
20865: waveform_sig_rx =986;
20866: waveform_sig_rx =827;
20867: waveform_sig_rx =756;
20868: waveform_sig_rx =980;
20869: waveform_sig_rx =933;
20870: waveform_sig_rx =739;
20871: waveform_sig_rx =890;
20872: waveform_sig_rx =1053;
20873: waveform_sig_rx =738;
20874: waveform_sig_rx =931;
20875: waveform_sig_rx =908;
20876: waveform_sig_rx =886;
20877: waveform_sig_rx =901;
20878: waveform_sig_rx =967;
20879: waveform_sig_rx =837;
20880: waveform_sig_rx =900;
20881: waveform_sig_rx =1126;
20882: waveform_sig_rx =681;
20883: waveform_sig_rx =1068;
20884: waveform_sig_rx =1046;
20885: waveform_sig_rx =718;
20886: waveform_sig_rx =1079;
20887: waveform_sig_rx =1068;
20888: waveform_sig_rx =721;
20889: waveform_sig_rx =1053;
20890: waveform_sig_rx =1075;
20891: waveform_sig_rx =800;
20892: waveform_sig_rx =1020;
20893: waveform_sig_rx =1040;
20894: waveform_sig_rx =984;
20895: waveform_sig_rx =808;
20896: waveform_sig_rx =1167;
20897: waveform_sig_rx =996;
20898: waveform_sig_rx =805;
20899: waveform_sig_rx =1106;
20900: waveform_sig_rx =1084;
20901: waveform_sig_rx =797;
20902: waveform_sig_rx =1095;
20903: waveform_sig_rx =1100;
20904: waveform_sig_rx =927;
20905: waveform_sig_rx =948;
20906: waveform_sig_rx =1148;
20907: waveform_sig_rx =1032;
20908: waveform_sig_rx =861;
20909: waveform_sig_rx =1153;
20910: waveform_sig_rx =1081;
20911: waveform_sig_rx =860;
20912: waveform_sig_rx =1094;
20913: waveform_sig_rx =1196;
20914: waveform_sig_rx =856;
20915: waveform_sig_rx =1144;
20916: waveform_sig_rx =1008;
20917: waveform_sig_rx =1046;
20918: waveform_sig_rx =1107;
20919: waveform_sig_rx =1098;
20920: waveform_sig_rx =984;
20921: waveform_sig_rx =1068;
20922: waveform_sig_rx =1219;
20923: waveform_sig_rx =835;
20924: waveform_sig_rx =1215;
20925: waveform_sig_rx =1115;
20926: waveform_sig_rx =908;
20927: waveform_sig_rx =1198;
20928: waveform_sig_rx =1187;
20929: waveform_sig_rx =902;
20930: waveform_sig_rx =1133;
20931: waveform_sig_rx =1240;
20932: waveform_sig_rx =924;
20933: waveform_sig_rx =1095;
20934: waveform_sig_rx =1247;
20935: waveform_sig_rx =1018;
20936: waveform_sig_rx =944;
20937: waveform_sig_rx =1339;
20938: waveform_sig_rx =1019;
20939: waveform_sig_rx =999;
20940: waveform_sig_rx =1214;
20941: waveform_sig_rx =1176;
20942: waveform_sig_rx =981;
20943: waveform_sig_rx =1155;
20944: waveform_sig_rx =1205;
20945: waveform_sig_rx =1034;
20946: waveform_sig_rx =1032;
20947: waveform_sig_rx =1286;
20948: waveform_sig_rx =1121;
20949: waveform_sig_rx =946;
20950: waveform_sig_rx =1291;
20951: waveform_sig_rx =1161;
20952: waveform_sig_rx =925;
20953: waveform_sig_rx =1225;
20954: waveform_sig_rx =1259;
20955: waveform_sig_rx =916;
20956: waveform_sig_rx =1276;
20957: waveform_sig_rx =1023;
20958: waveform_sig_rx =1164;
20959: waveform_sig_rx =1165;
20960: waveform_sig_rx =1119;
20961: waveform_sig_rx =1108;
20962: waveform_sig_rx =1119;
20963: waveform_sig_rx =1267;
20964: waveform_sig_rx =953;
20965: waveform_sig_rx =1258;
20966: waveform_sig_rx =1220;
20967: waveform_sig_rx =970;
20968: waveform_sig_rx =1231;
20969: waveform_sig_rx =1276;
20970: waveform_sig_rx =903;
20971: waveform_sig_rx =1214;
20972: waveform_sig_rx =1302;
20973: waveform_sig_rx =919;
20974: waveform_sig_rx =1207;
20975: waveform_sig_rx =1292;
20976: waveform_sig_rx =1034;
20977: waveform_sig_rx =1048;
20978: waveform_sig_rx =1356;
20979: waveform_sig_rx =1042;
20980: waveform_sig_rx =1085;
20981: waveform_sig_rx =1211;
20982: waveform_sig_rx =1228;
20983: waveform_sig_rx =1020;
20984: waveform_sig_rx =1168;
20985: waveform_sig_rx =1264;
20986: waveform_sig_rx =1049;
20987: waveform_sig_rx =1049;
20988: waveform_sig_rx =1342;
20989: waveform_sig_rx =1095;
20990: waveform_sig_rx =971;
20991: waveform_sig_rx =1365;
20992: waveform_sig_rx =1106;
20993: waveform_sig_rx =977;
20994: waveform_sig_rx =1278;
20995: waveform_sig_rx =1174;
20996: waveform_sig_rx =1004;
20997: waveform_sig_rx =1264;
20998: waveform_sig_rx =1000;
20999: waveform_sig_rx =1253;
21000: waveform_sig_rx =1078;
21001: waveform_sig_rx =1180;
21002: waveform_sig_rx =1108;
21003: waveform_sig_rx =1082;
21004: waveform_sig_rx =1322;
21005: waveform_sig_rx =900;
21006: waveform_sig_rx =1231;
21007: waveform_sig_rx =1242;
21008: waveform_sig_rx =881;
21009: waveform_sig_rx =1277;
21010: waveform_sig_rx =1223;
21011: waveform_sig_rx =881;
21012: waveform_sig_rx =1248;
21013: waveform_sig_rx =1255;
21014: waveform_sig_rx =913;
21015: waveform_sig_rx =1188;
21016: waveform_sig_rx =1291;
21017: waveform_sig_rx =964;
21018: waveform_sig_rx =1081;
21019: waveform_sig_rx =1287;
21020: waveform_sig_rx =1017;
21021: waveform_sig_rx =1100;
21022: waveform_sig_rx =1095;
21023: waveform_sig_rx =1242;
21024: waveform_sig_rx =950;
21025: waveform_sig_rx =1093;
21026: waveform_sig_rx =1312;
21027: waveform_sig_rx =933;
21028: waveform_sig_rx =1081;
21029: waveform_sig_rx =1313;
21030: waveform_sig_rx =972;
21031: waveform_sig_rx =1020;
21032: waveform_sig_rx =1249;
21033: waveform_sig_rx =1049;
21034: waveform_sig_rx =987;
21035: waveform_sig_rx =1158;
21036: waveform_sig_rx =1156;
21037: waveform_sig_rx =936;
21038: waveform_sig_rx =1153;
21039: waveform_sig_rx =974;
21040: waveform_sig_rx =1167;
21041: waveform_sig_rx =986;
21042: waveform_sig_rx =1152;
21043: waveform_sig_rx =987;
21044: waveform_sig_rx =1048;
21045: waveform_sig_rx =1263;
21046: waveform_sig_rx =783;
21047: waveform_sig_rx =1229;
21048: waveform_sig_rx =1133;
21049: waveform_sig_rx =766;
21050: waveform_sig_rx =1249;
21051: waveform_sig_rx =1107;
21052: waveform_sig_rx =778;
21053: waveform_sig_rx =1199;
21054: waveform_sig_rx =1087;
21055: waveform_sig_rx =828;
21056: waveform_sig_rx =1131;
21057: waveform_sig_rx =1092;
21058: waveform_sig_rx =900;
21059: waveform_sig_rx =974;
21060: waveform_sig_rx =1151;
21061: waveform_sig_rx =960;
21062: waveform_sig_rx =915;
21063: waveform_sig_rx =1018;
21064: waveform_sig_rx =1159;
21065: waveform_sig_rx =751;
21066: waveform_sig_rx =1073;
21067: waveform_sig_rx =1133;
21068: waveform_sig_rx =768;
21069: waveform_sig_rx =1036;
21070: waveform_sig_rx =1107;
21071: waveform_sig_rx =865;
21072: waveform_sig_rx =913;
21073: waveform_sig_rx =1057;
21074: waveform_sig_rx =980;
21075: waveform_sig_rx =811;
21076: waveform_sig_rx =1027;
21077: waveform_sig_rx =1053;
21078: waveform_sig_rx =787;
21079: waveform_sig_rx =1045;
21080: waveform_sig_rx =852;
21081: waveform_sig_rx =1007;
21082: waveform_sig_rx =872;
21083: waveform_sig_rx =1041;
21084: waveform_sig_rx =803;
21085: waveform_sig_rx =952;
21086: waveform_sig_rx =1074;
21087: waveform_sig_rx =616;
21088: waveform_sig_rx =1110;
21089: waveform_sig_rx =920;
21090: waveform_sig_rx =641;
21091: waveform_sig_rx =1149;
21092: waveform_sig_rx =867;
21093: waveform_sig_rx =682;
21094: waveform_sig_rx =1055;
21095: waveform_sig_rx =870;
21096: waveform_sig_rx =753;
21097: waveform_sig_rx =903;
21098: waveform_sig_rx =956;
21099: waveform_sig_rx =764;
21100: waveform_sig_rx =743;
21101: waveform_sig_rx =1037;
21102: waveform_sig_rx =767;
21103: waveform_sig_rx =747;
21104: waveform_sig_rx =934;
21105: waveform_sig_rx =912;
21106: waveform_sig_rx =610;
21107: waveform_sig_rx =942;
21108: waveform_sig_rx =904;
21109: waveform_sig_rx =639;
21110: waveform_sig_rx =837;
21111: waveform_sig_rx =894;
21112: waveform_sig_rx =707;
21113: waveform_sig_rx =693;
21114: waveform_sig_rx =908;
21115: waveform_sig_rx =788;
21116: waveform_sig_rx =597;
21117: waveform_sig_rx =879;
21118: waveform_sig_rx =859;
21119: waveform_sig_rx =556;
21120: waveform_sig_rx =879;
21121: waveform_sig_rx =636;
21122: waveform_sig_rx =769;
21123: waveform_sig_rx =698;
21124: waveform_sig_rx =782;
21125: waveform_sig_rx =583;
21126: waveform_sig_rx =800;
21127: waveform_sig_rx =776;
21128: waveform_sig_rx =462;
21129: waveform_sig_rx =901;
21130: waveform_sig_rx =643;
21131: waveform_sig_rx =513;
21132: waveform_sig_rx =871;
21133: waveform_sig_rx =644;
21134: waveform_sig_rx =502;
21135: waveform_sig_rx =777;
21136: waveform_sig_rx =681;
21137: waveform_sig_rx =525;
21138: waveform_sig_rx =656;
21139: waveform_sig_rx =767;
21140: waveform_sig_rx =480;
21141: waveform_sig_rx =526;
21142: waveform_sig_rx =826;
21143: waveform_sig_rx =461;
21144: waveform_sig_rx =529;
21145: waveform_sig_rx =703;
21146: waveform_sig_rx =612;
21147: waveform_sig_rx =428;
21148: waveform_sig_rx =694;
21149: waveform_sig_rx =618;
21150: waveform_sig_rx =447;
21151: waveform_sig_rx =544;
21152: waveform_sig_rx =671;
21153: waveform_sig_rx =476;
21154: waveform_sig_rx =415;
21155: waveform_sig_rx =707;
21156: waveform_sig_rx =508;
21157: waveform_sig_rx =321;
21158: waveform_sig_rx =667;
21159: waveform_sig_rx =539;
21160: waveform_sig_rx =327;
21161: waveform_sig_rx =649;
21162: waveform_sig_rx =350;
21163: waveform_sig_rx =553;
21164: waveform_sig_rx =435;
21165: waveform_sig_rx =507;
21166: waveform_sig_rx =344;
21167: waveform_sig_rx =544;
21168: waveform_sig_rx =471;
21169: waveform_sig_rx =248;
21170: waveform_sig_rx =628;
21171: waveform_sig_rx =385;
21172: waveform_sig_rx =286;
21173: waveform_sig_rx =542;
21174: waveform_sig_rx =416;
21175: waveform_sig_rx =217;
21176: waveform_sig_rx =493;
21177: waveform_sig_rx =477;
21178: waveform_sig_rx =170;
21179: waveform_sig_rx =441;
21180: waveform_sig_rx =522;
21181: waveform_sig_rx =143;
21182: waveform_sig_rx =332;
21183: waveform_sig_rx =521;
21184: waveform_sig_rx =180;
21185: waveform_sig_rx =287;
21186: waveform_sig_rx =386;
21187: waveform_sig_rx =344;
21188: waveform_sig_rx =151;
21189: waveform_sig_rx =367;
21190: waveform_sig_rx =372;
21191: waveform_sig_rx =142;
21192: waveform_sig_rx =250;
21193: waveform_sig_rx =450;
21194: waveform_sig_rx =154;
21195: waveform_sig_rx =133;
21196: waveform_sig_rx =446;
21197: waveform_sig_rx =164;
21198: waveform_sig_rx =68;
21199: waveform_sig_rx =400;
21200: waveform_sig_rx =199;
21201: waveform_sig_rx =81;
21202: waveform_sig_rx =323;
21203: waveform_sig_rx =23;
21204: waveform_sig_rx =319;
21205: waveform_sig_rx =102;
21206: waveform_sig_rx =231;
21207: waveform_sig_rx =53;
21208: waveform_sig_rx =203;
21209: waveform_sig_rx =200;
21210: waveform_sig_rx =-49;
21211: waveform_sig_rx =273;
21212: waveform_sig_rx =127;
21213: waveform_sig_rx =-59;
21214: waveform_sig_rx =244;
21215: waveform_sig_rx =174;
21216: waveform_sig_rx =-165;
21217: waveform_sig_rx =274;
21218: waveform_sig_rx =147;
21219: waveform_sig_rx =-169;
21220: waveform_sig_rx =233;
21221: waveform_sig_rx =115;
21222: waveform_sig_rx =-133;
21223: waveform_sig_rx =85;
21224: waveform_sig_rx =136;
21225: waveform_sig_rx =-55;
21226: waveform_sig_rx =-16;
21227: waveform_sig_rx =74;
21228: waveform_sig_rx =64;
21229: waveform_sig_rx =-198;
21230: waveform_sig_rx =90;
21231: waveform_sig_rx =81;
21232: waveform_sig_rx =-171;
21233: waveform_sig_rx =-35;
21234: waveform_sig_rx =129;
21235: waveform_sig_rx =-193;
21236: waveform_sig_rx =-162;
21237: waveform_sig_rx =157;
21238: waveform_sig_rx =-202;
21239: waveform_sig_rx =-182;
21240: waveform_sig_rx =78;
21241: waveform_sig_rx =-150;
21242: waveform_sig_rx =-158;
21243: waveform_sig_rx =-65;
21244: waveform_sig_rx =-222;
21245: waveform_sig_rx =24;
21246: waveform_sig_rx =-276;
21247: waveform_sig_rx =-1;
21248: waveform_sig_rx =-283;
21249: waveform_sig_rx =-109;
21250: waveform_sig_rx =-60;
21251: waveform_sig_rx =-406;
21252: waveform_sig_rx =9;
21253: waveform_sig_rx =-166;
21254: waveform_sig_rx =-433;
21255: waveform_sig_rx =78;
21256: waveform_sig_rx =-212;
21257: waveform_sig_rx =-451;
21258: waveform_sig_rx =42;
21259: waveform_sig_rx =-244;
21260: waveform_sig_rx =-418;
21261: waveform_sig_rx =-103;
21262: waveform_sig_rx =-213;
21263: waveform_sig_rx =-405;
21264: waveform_sig_rx =-257;
21265: waveform_sig_rx =-147;
21266: waveform_sig_rx =-367;
21267: waveform_sig_rx =-355;
21268: waveform_sig_rx =-209;
21269: waveform_sig_rx =-263;
21270: waveform_sig_rx =-495;
21271: waveform_sig_rx =-211;
21272: waveform_sig_rx =-224;
21273: waveform_sig_rx =-539;
21274: waveform_sig_rx =-296;
21275: waveform_sig_rx =-163;
21276: waveform_sig_rx =-584;
21277: waveform_sig_rx =-347;
21278: waveform_sig_rx =-236;
21279: waveform_sig_rx =-495;
21280: waveform_sig_rx =-425;
21281: waveform_sig_rx =-341;
21282: waveform_sig_rx =-348;
21283: waveform_sig_rx =-515;
21284: waveform_sig_rx =-388;
21285: waveform_sig_rx =-441;
21286: waveform_sig_rx =-402;
21287: waveform_sig_rx =-525;
21288: waveform_sig_rx =-293;
21289: waveform_sig_rx =-672;
21290: waveform_sig_rx =-290;
21291: waveform_sig_rx =-425;
21292: waveform_sig_rx =-696;
21293: waveform_sig_rx =-222;
21294: waveform_sig_rx =-571;
21295: waveform_sig_rx =-647;
21296: waveform_sig_rx =-276;
21297: waveform_sig_rx =-557;
21298: waveform_sig_rx =-708;
21299: waveform_sig_rx =-296;
21300: waveform_sig_rx =-553;
21301: waveform_sig_rx =-687;
21302: waveform_sig_rx =-391;
21303: waveform_sig_rx =-528;
21304: waveform_sig_rx =-667;
21305: waveform_sig_rx =-547;
21306: waveform_sig_rx =-444;
21307: waveform_sig_rx =-615;
21308: waveform_sig_rx =-682;
21309: waveform_sig_rx =-431;
21310: waveform_sig_rx =-542;
21311: waveform_sig_rx =-818;
21312: waveform_sig_rx =-390;
21313: waveform_sig_rx =-593;
21314: waveform_sig_rx =-799;
21315: waveform_sig_rx =-510;
21316: waveform_sig_rx =-549;
21317: waveform_sig_rx =-742;
21318: waveform_sig_rx =-644;
21319: waveform_sig_rx =-518;
21320: waveform_sig_rx =-680;
21321: waveform_sig_rx =-784;
21322: waveform_sig_rx =-541;
21323: waveform_sig_rx =-599;
21324: waveform_sig_rx =-841;
21325: waveform_sig_rx =-555;
21326: waveform_sig_rx =-774;
21327: waveform_sig_rx =-662;
21328: waveform_sig_rx =-701;
21329: waveform_sig_rx =-627;
21330: waveform_sig_rx =-898;
21331: waveform_sig_rx =-527;
21332: waveform_sig_rx =-778;
21333: waveform_sig_rx =-889;
21334: waveform_sig_rx =-506;
21335: waveform_sig_rx =-855;
21336: waveform_sig_rx =-878;
21337: waveform_sig_rx =-531;
21338: waveform_sig_rx =-821;
21339: waveform_sig_rx =-950;
21340: waveform_sig_rx =-551;
21341: waveform_sig_rx =-857;
21342: waveform_sig_rx =-884;
21343: waveform_sig_rx =-684;
21344: waveform_sig_rx =-758;
21345: waveform_sig_rx =-900;
21346: waveform_sig_rx =-864;
21347: waveform_sig_rx =-611;
21348: waveform_sig_rx =-941;
21349: waveform_sig_rx =-933;
21350: waveform_sig_rx =-589;
21351: waveform_sig_rx =-918;
21352: waveform_sig_rx =-974;
21353: waveform_sig_rx =-658;
21354: waveform_sig_rx =-902;
21355: waveform_sig_rx =-924;
21356: waveform_sig_rx =-849;
21357: waveform_sig_rx =-721;
21358: waveform_sig_rx =-977;
21359: waveform_sig_rx =-957;
21360: waveform_sig_rx =-661;
21361: waveform_sig_rx =-983;
21362: waveform_sig_rx =-999;
21363: waveform_sig_rx =-700;
21364: waveform_sig_rx =-909;
21365: waveform_sig_rx =-1011;
21366: waveform_sig_rx =-801;
21367: waveform_sig_rx =-1005;
21368: waveform_sig_rx =-864;
21369: waveform_sig_rx =-947;
21370: waveform_sig_rx =-865;
21371: waveform_sig_rx =-1113;
21372: waveform_sig_rx =-752;
21373: waveform_sig_rx =-1018;
21374: waveform_sig_rx =-1074;
21375: waveform_sig_rx =-742;
21376: waveform_sig_rx =-1087;
21377: waveform_sig_rx =-1021;
21378: waveform_sig_rx =-796;
21379: waveform_sig_rx =-1011;
21380: waveform_sig_rx =-1115;
21381: waveform_sig_rx =-826;
21382: waveform_sig_rx =-984;
21383: waveform_sig_rx =-1154;
21384: waveform_sig_rx =-889;
21385: waveform_sig_rx =-888;
21386: waveform_sig_rx =-1227;
21387: waveform_sig_rx =-960;
21388: waveform_sig_rx =-846;
21389: waveform_sig_rx =-1178;
21390: waveform_sig_rx =-1025;
21391: waveform_sig_rx =-881;
21392: waveform_sig_rx =-1069;
21393: waveform_sig_rx =-1110;
21394: waveform_sig_rx =-913;
21395: waveform_sig_rx =-1001;
21396: waveform_sig_rx =-1158;
21397: waveform_sig_rx =-1025;
21398: waveform_sig_rx =-890;
21399: waveform_sig_rx =-1230;
21400: waveform_sig_rx =-1095;
21401: waveform_sig_rx =-844;
21402: waveform_sig_rx =-1211;
21403: waveform_sig_rx =-1158;
21404: waveform_sig_rx =-885;
21405: waveform_sig_rx =-1120;
21406: waveform_sig_rx =-1146;
21407: waveform_sig_rx =-984;
21408: waveform_sig_rx =-1203;
21409: waveform_sig_rx =-974;
21410: waveform_sig_rx =-1159;
21411: waveform_sig_rx =-1033;
21412: waveform_sig_rx =-1228;
21413: waveform_sig_rx =-949;
21414: waveform_sig_rx =-1145;
21415: waveform_sig_rx =-1214;
21416: waveform_sig_rx =-932;
21417: waveform_sig_rx =-1181;
21418: waveform_sig_rx =-1218;
21419: waveform_sig_rx =-930;
21420: waveform_sig_rx =-1121;
21421: waveform_sig_rx =-1311;
21422: waveform_sig_rx =-871;
21423: waveform_sig_rx =-1148;
21424: waveform_sig_rx =-1301;
21425: waveform_sig_rx =-948;
21426: waveform_sig_rx =-1103;
21427: waveform_sig_rx =-1318;
21428: waveform_sig_rx =-1016;
21429: waveform_sig_rx =-1065;
21430: waveform_sig_rx =-1256;
21431: waveform_sig_rx =-1170;
21432: waveform_sig_rx =-1046;
21433: waveform_sig_rx =-1146;
21434: waveform_sig_rx =-1287;
21435: waveform_sig_rx =-1013;
21436: waveform_sig_rx =-1107;
21437: waveform_sig_rx =-1306;
21438: waveform_sig_rx =-1071;
21439: waveform_sig_rx =-997;
21440: waveform_sig_rx =-1332;
21441: waveform_sig_rx =-1144;
21442: waveform_sig_rx =-980;
21443: waveform_sig_rx =-1314;
21444: waveform_sig_rx =-1195;
21445: waveform_sig_rx =-987;
21446: waveform_sig_rx =-1231;
21447: waveform_sig_rx =-1182;
21448: waveform_sig_rx =-1117;
21449: waveform_sig_rx =-1252;
21450: waveform_sig_rx =-1029;
21451: waveform_sig_rx =-1275;
21452: waveform_sig_rx =-1037;
21453: waveform_sig_rx =-1334;
21454: waveform_sig_rx =-1023;
21455: waveform_sig_rx =-1178;
21456: waveform_sig_rx =-1319;
21457: waveform_sig_rx =-947;
21458: waveform_sig_rx =-1253;
21459: waveform_sig_rx =-1305;
21460: waveform_sig_rx =-891;
21461: waveform_sig_rx =-1254;
21462: waveform_sig_rx =-1321;
21463: waveform_sig_rx =-891;
21464: waveform_sig_rx =-1278;
21465: waveform_sig_rx =-1280;
21466: waveform_sig_rx =-977;
21467: waveform_sig_rx =-1144;
21468: waveform_sig_rx =-1323;
21469: waveform_sig_rx =-1054;
21470: waveform_sig_rx =-1101;
21471: waveform_sig_rx =-1246;
21472: waveform_sig_rx =-1206;
21473: waveform_sig_rx =-1054;
21474: waveform_sig_rx =-1145;
21475: waveform_sig_rx =-1336;
21476: waveform_sig_rx =-987;
21477: waveform_sig_rx =-1129;
21478: waveform_sig_rx =-1351;
21479: waveform_sig_rx =-1020;
21480: waveform_sig_rx =-1071;
21481: waveform_sig_rx =-1343;
21482: waveform_sig_rx =-1074;
21483: waveform_sig_rx =-1056;
21484: waveform_sig_rx =-1250;
21485: waveform_sig_rx =-1180;
21486: waveform_sig_rx =-1032;
21487: waveform_sig_rx =-1191;
21488: waveform_sig_rx =-1228;
21489: waveform_sig_rx =-1111;
21490: waveform_sig_rx =-1205;
21491: waveform_sig_rx =-1073;
21492: waveform_sig_rx =-1214;
21493: waveform_sig_rx =-1024;
21494: waveform_sig_rx =-1319;
21495: waveform_sig_rx =-942;
21496: waveform_sig_rx =-1200;
21497: waveform_sig_rx =-1301;
21498: waveform_sig_rx =-882;
21499: waveform_sig_rx =-1284;
21500: waveform_sig_rx =-1245;
21501: waveform_sig_rx =-853;
21502: waveform_sig_rx =-1316;
21503: waveform_sig_rx =-1223;
21504: waveform_sig_rx =-883;
21505: waveform_sig_rx =-1266;
21506: waveform_sig_rx =-1161;
21507: waveform_sig_rx =-1010;
21508: waveform_sig_rx =-1099;
21509: waveform_sig_rx =-1258;
21510: waveform_sig_rx =-1051;
21511: waveform_sig_rx =-1026;
21512: waveform_sig_rx =-1218;
21513: waveform_sig_rx =-1169;
21514: waveform_sig_rx =-950;
21515: waveform_sig_rx =-1144;
21516: waveform_sig_rx =-1261;
21517: waveform_sig_rx =-896;
21518: waveform_sig_rx =-1137;
21519: waveform_sig_rx =-1245;
21520: waveform_sig_rx =-964;
21521: waveform_sig_rx =-1073;
21522: waveform_sig_rx =-1210;
21523: waveform_sig_rx =-1055;
21524: waveform_sig_rx =-983;
21525: waveform_sig_rx =-1166;
21526: waveform_sig_rx =-1157;
21527: waveform_sig_rx =-900;
21528: waveform_sig_rx =-1123;
21529: waveform_sig_rx =-1144;
21530: waveform_sig_rx =-997;
21531: waveform_sig_rx =-1123;
21532: waveform_sig_rx =-1016;
21533: waveform_sig_rx =-1077;
21534: waveform_sig_rx =-982;
21535: waveform_sig_rx =-1245;
21536: waveform_sig_rx =-790;
21537: waveform_sig_rx =-1182;
21538: waveform_sig_rx =-1143;
21539: waveform_sig_rx =-775;
21540: waveform_sig_rx =-1246;
21541: waveform_sig_rx =-1049;
21542: waveform_sig_rx =-814;
21543: waveform_sig_rx =-1207;
21544: waveform_sig_rx =-1057;
21545: waveform_sig_rx =-836;
21546: waveform_sig_rx =-1102;
21547: waveform_sig_rx =-1065;
21548: waveform_sig_rx =-917;
21549: waveform_sig_rx =-935;
21550: waveform_sig_rx =-1207;
21551: waveform_sig_rx =-890;
21552: waveform_sig_rx =-881;
21553: waveform_sig_rx =-1115;
21554: waveform_sig_rx =-985;
21555: waveform_sig_rx =-811;
21556: waveform_sig_rx =-1058;
21557: waveform_sig_rx =-1081;
21558: waveform_sig_rx =-762;
21559: waveform_sig_rx =-1024;
21560: waveform_sig_rx =-1053;
21561: waveform_sig_rx =-823;
21562: waveform_sig_rx =-919;
21563: waveform_sig_rx =-1042;
21564: waveform_sig_rx =-924;
21565: waveform_sig_rx =-782;
21566: waveform_sig_rx =-1026;
21567: waveform_sig_rx =-1043;
21568: waveform_sig_rx =-684;
21569: waveform_sig_rx =-1028;
21570: waveform_sig_rx =-957;
21571: waveform_sig_rx =-821;
21572: waveform_sig_rx =-1018;
21573: waveform_sig_rx =-809;
21574: waveform_sig_rx =-916;
21575: waveform_sig_rx =-866;
21576: waveform_sig_rx =-1037;
21577: waveform_sig_rx =-652;
21578: waveform_sig_rx =-1059;
21579: waveform_sig_rx =-877;
21580: waveform_sig_rx =-684;
21581: waveform_sig_rx =-1072;
21582: waveform_sig_rx =-827;
21583: waveform_sig_rx =-694;
21584: waveform_sig_rx =-961;
21585: waveform_sig_rx =-899;
21586: waveform_sig_rx =-672;
21587: waveform_sig_rx =-889;
21588: waveform_sig_rx =-918;
21589: waveform_sig_rx =-699;
21590: waveform_sig_rx =-764;
21591: waveform_sig_rx =-1035;
21592: waveform_sig_rx =-647;
21593: waveform_sig_rx =-737;
21594: waveform_sig_rx =-936;
21595: waveform_sig_rx =-776;
21596: waveform_sig_rx =-647;
21597: waveform_sig_rx =-866;
21598: waveform_sig_rx =-821;
21599: waveform_sig_rx =-612;
21600: waveform_sig_rx =-818;
21601: waveform_sig_rx =-844;
21602: waveform_sig_rx =-662;
21603: waveform_sig_rx =-661;
21604: waveform_sig_rx =-880;
21605: waveform_sig_rx =-719;
21606: waveform_sig_rx =-512;
21607: waveform_sig_rx =-882;
21608: waveform_sig_rx =-769;
21609: waveform_sig_rx =-468;
21610: waveform_sig_rx =-894;
21611: waveform_sig_rx =-645;
21612: waveform_sig_rx =-652;
21613: waveform_sig_rx =-793;
21614: waveform_sig_rx =-562;
21615: waveform_sig_rx =-765;
21616: waveform_sig_rx =-614;
21617: waveform_sig_rx =-800;
21618: waveform_sig_rx =-487;
21619: waveform_sig_rx =-797;
21620: waveform_sig_rx =-672;
21621: waveform_sig_rx =-474;
21622: waveform_sig_rx =-795;
21623: waveform_sig_rx =-644;
21624: waveform_sig_rx =-449;
21625: waveform_sig_rx =-729;
21626: waveform_sig_rx =-683;
21627: waveform_sig_rx =-423;
21628: waveform_sig_rx =-675;
21629: waveform_sig_rx =-708;
21630: waveform_sig_rx =-410;
21631: waveform_sig_rx =-552;
21632: waveform_sig_rx =-812;
21633: waveform_sig_rx =-355;
21634: waveform_sig_rx =-559;
21635: waveform_sig_rx =-652;
21636: waveform_sig_rx =-503;
21637: waveform_sig_rx =-462;
21638: waveform_sig_rx =-570;
21639: waveform_sig_rx =-608;
21640: waveform_sig_rx =-382;
21641: waveform_sig_rx =-528;
21642: waveform_sig_rx =-660;
21643: waveform_sig_rx =-363;
21644: waveform_sig_rx =-409;
21645: waveform_sig_rx =-692;
21646: waveform_sig_rx =-402;
21647: waveform_sig_rx =-354;
21648: waveform_sig_rx =-649;
21649: waveform_sig_rx =-458;
21650: waveform_sig_rx =-280;
21651: waveform_sig_rx =-596;
21652: waveform_sig_rx =-385;
21653: waveform_sig_rx =-456;
21654: waveform_sig_rx =-488;
21655: waveform_sig_rx =-321;
21656: waveform_sig_rx =-501;
21657: waveform_sig_rx =-325;
21658: waveform_sig_rx =-543;
21659: waveform_sig_rx =-191;
21660: waveform_sig_rx =-502;
21661: waveform_sig_rx =-421;
21662: waveform_sig_rx =-167;
21663: waveform_sig_rx =-517;
21664: waveform_sig_rx =-410;
21665: waveform_sig_rx =-118;
21666: waveform_sig_rx =-506;
21667: waveform_sig_rx =-444;
21668: waveform_sig_rx =-71;
21669: waveform_sig_rx =-500;
21670: waveform_sig_rx =-386;
21671: waveform_sig_rx =-123;
21672: waveform_sig_rx =-365;
21673: waveform_sig_rx =-437;
21674: waveform_sig_rx =-113;
21675: waveform_sig_rx =-279;
21676: waveform_sig_rx =-341;
21677: waveform_sig_rx =-278;
21678: waveform_sig_rx =-125;
21679: waveform_sig_rx =-295;
21680: waveform_sig_rx =-353;
21681: waveform_sig_rx =-40;
21682: waveform_sig_rx =-269;
21683: waveform_sig_rx =-388;
21684: waveform_sig_rx =-56;
21685: waveform_sig_rx =-174;
21686: waveform_sig_rx =-396;
21687: waveform_sig_rx =-90;
21688: waveform_sig_rx =-104;
21689: waveform_sig_rx =-342;
21690: waveform_sig_rx =-138;
21691: waveform_sig_rx =-25;
21692: waveform_sig_rx =-279;
21693: waveform_sig_rx =-119;
21694: waveform_sig_rx =-171;
21695: waveform_sig_rx =-126;
21696: waveform_sig_rx =-109;
21697: waveform_sig_rx =-169;
21698: waveform_sig_rx =-16;
21699: waveform_sig_rx =-302;
21700: waveform_sig_rx =120;
21701: waveform_sig_rx =-245;
21702: waveform_sig_rx =-144;
21703: waveform_sig_rx =158;
21704: waveform_sig_rx =-273;
21705: waveform_sig_rx =-72;
21706: waveform_sig_rx =186;
21707: waveform_sig_rx =-294;
21708: waveform_sig_rx =-45;
21709: waveform_sig_rx =212;
21710: waveform_sig_rx =-211;
21711: waveform_sig_rx =-2;
21712: waveform_sig_rx =116;
21713: waveform_sig_rx =-31;
21714: waveform_sig_rx =-114;
21715: waveform_sig_rx =119;
21716: waveform_sig_rx =53;
21717: waveform_sig_rx =-80;
21718: waveform_sig_rx =-1;
21719: waveform_sig_rx =200;
21720: waveform_sig_rx =-73;
21721: waveform_sig_rx =-19;
21722: waveform_sig_rx =251;
21723: waveform_sig_rx =-24;
21724: waveform_sig_rx =-78;
21725: waveform_sig_rx =254;
21726: waveform_sig_rx =79;
21727: waveform_sig_rx =-95;
21728: waveform_sig_rx =219;
21729: waveform_sig_rx =141;
21730: waveform_sig_rx =4;
21731: waveform_sig_rx =120;
21732: waveform_sig_rx =252;
21733: waveform_sig_rx =90;
21734: waveform_sig_rx =118;
21735: waveform_sig_rx =183;
21736: waveform_sig_rx =185;
21737: waveform_sig_rx =124;
21738: waveform_sig_rx =215;
21739: waveform_sig_rx =184;
21740: waveform_sig_rx =30;
21741: waveform_sig_rx =463;
21742: waveform_sig_rx =-36;
21743: waveform_sig_rx =227;
21744: waveform_sig_rx =390;
21745: waveform_sig_rx =-14;
21746: waveform_sig_rx =286;
21747: waveform_sig_rx =404;
21748: waveform_sig_rx =52;
21749: waveform_sig_rx =249;
21750: waveform_sig_rx =473;
21751: waveform_sig_rx =80;
21752: waveform_sig_rx =272;
21753: waveform_sig_rx =395;
21754: waveform_sig_rx =245;
21755: waveform_sig_rx =176;
21756: waveform_sig_rx =403;
21757: waveform_sig_rx =343;
21758: waveform_sig_rx =216;
21759: waveform_sig_rx =292;
21760: waveform_sig_rx =552;
21761: waveform_sig_rx =155;
21762: waveform_sig_rx =323;
21763: waveform_sig_rx =575;
21764: waveform_sig_rx =195;
21765: waveform_sig_rx =321;
21766: waveform_sig_rx =493;
21767: waveform_sig_rx =377;
21768: waveform_sig_rx =273;
21769: waveform_sig_rx =454;
21770: waveform_sig_rx =507;
21771: waveform_sig_rx =269;
21772: waveform_sig_rx =366;
21773: waveform_sig_rx =618;
21774: waveform_sig_rx =280;
21775: waveform_sig_rx =433;
21776: waveform_sig_rx =483;
21777: waveform_sig_rx =403;
21778: waveform_sig_rx =488;
21779: waveform_sig_rx =497;
21780: waveform_sig_rx =428;
21781: waveform_sig_rx =398;
21782: waveform_sig_rx =697;
21783: waveform_sig_rx =249;
21784: waveform_sig_rx =568;
21785: waveform_sig_rx =635;
21786: waveform_sig_rx =289;
21787: waveform_sig_rx =572;
21788: waveform_sig_rx =684;
21789: waveform_sig_rx =328;
21790: waveform_sig_rx =541;
21791: waveform_sig_rx =719;
21792: waveform_sig_rx =361;
21793: waveform_sig_rx =547;
21794: waveform_sig_rx =637;
21795: waveform_sig_rx =558;
21796: waveform_sig_rx =393;
21797: waveform_sig_rx =715;
21798: waveform_sig_rx =656;
21799: waveform_sig_rx =385;
21800: waveform_sig_rx =648;
21801: waveform_sig_rx =767;
21802: waveform_sig_rx =386;
21803: waveform_sig_rx =674;
21804: waveform_sig_rx =714;
21805: waveform_sig_rx =523;
21806: waveform_sig_rx =576;
21807: waveform_sig_rx =706;
21808: waveform_sig_rx =719;
21809: waveform_sig_rx =455;
21810: waveform_sig_rx =746;
21811: waveform_sig_rx =795;
21812: waveform_sig_rx =440;
21813: waveform_sig_rx =713;
21814: waveform_sig_rx =829;
21815: waveform_sig_rx =482;
21816: waveform_sig_rx =725;
21817: waveform_sig_rx =663;
21818: waveform_sig_rx =666;
21819: waveform_sig_rx =734;
21820: waveform_sig_rx =712;
21821: waveform_sig_rx =663;
21822: waveform_sig_rx =668;
21823: waveform_sig_rx =900;
21824: waveform_sig_rx =517;
21825: waveform_sig_rx =819;
21826: waveform_sig_rx =838;
21827: waveform_sig_rx =571;
21828: waveform_sig_rx =815;
21829: waveform_sig_rx =878;
21830: waveform_sig_rx =609;
21831: waveform_sig_rx =749;
21832: waveform_sig_rx =944;
21833: waveform_sig_rx =631;
21834: waveform_sig_rx =742;
21835: waveform_sig_rx =959;
21836: waveform_sig_rx =771;
21837: waveform_sig_rx =611;
21838: waveform_sig_rx =1036;
21839: waveform_sig_rx =780;
21840: waveform_sig_rx =682;
21841: waveform_sig_rx =910;
21842: waveform_sig_rx =892;
21843: waveform_sig_rx =722;
21844: waveform_sig_rx =848;
21845: waveform_sig_rx =944;
21846: waveform_sig_rx =828;
21847: waveform_sig_rx =741;
21848: waveform_sig_rx =1024;
21849: waveform_sig_rx =905;
21850: waveform_sig_rx =659;
21851: waveform_sig_rx =1024;
21852: waveform_sig_rx =932;
21853: waveform_sig_rx =704;
21854: waveform_sig_rx =945;
21855: waveform_sig_rx =1048;
21856: waveform_sig_rx =728;
21857: waveform_sig_rx =975;
21858: waveform_sig_rx =873;
21859: waveform_sig_rx =882;
21860: waveform_sig_rx =968;
21861: waveform_sig_rx =905;
21862: waveform_sig_rx =896;
21863: waveform_sig_rx =891;
21864: waveform_sig_rx =1075;
21865: waveform_sig_rx =769;
21866: waveform_sig_rx =998;
21867: waveform_sig_rx =1030;
21868: waveform_sig_rx =826;
21869: waveform_sig_rx =973;
21870: waveform_sig_rx =1162;
21871: waveform_sig_rx =778;
21872: waveform_sig_rx =934;
21873: waveform_sig_rx =1232;
21874: waveform_sig_rx =726;
21875: waveform_sig_rx =997;
21876: waveform_sig_rx =1163;
21877: waveform_sig_rx =855;
21878: waveform_sig_rx =882;
21879: waveform_sig_rx =1159;
21880: waveform_sig_rx =930;
21881: waveform_sig_rx =931;
21882: waveform_sig_rx =1028;
21883: waveform_sig_rx =1113;
21884: waveform_sig_rx =885;
21885: waveform_sig_rx =988;
21886: waveform_sig_rx =1176;
21887: waveform_sig_rx =948;
21888: waveform_sig_rx =889;
21889: waveform_sig_rx =1206;
21890: waveform_sig_rx =1020;
21891: waveform_sig_rx =823;
21892: waveform_sig_rx =1225;
21893: waveform_sig_rx =1055;
21894: waveform_sig_rx =874;
21895: waveform_sig_rx =1125;
21896: waveform_sig_rx =1139;
21897: waveform_sig_rx =916;
21898: waveform_sig_rx =1148;
21899: waveform_sig_rx =960;
21900: waveform_sig_rx =1119;
21901: waveform_sig_rx =1057;
21902: waveform_sig_rx =1063;
21903: waveform_sig_rx =1087;
21904: waveform_sig_rx =975;
21905: waveform_sig_rx =1268;
21906: waveform_sig_rx =886;
21907: waveform_sig_rx =1099;
21908: waveform_sig_rx =1237;
21909: waveform_sig_rx =861;
21910: waveform_sig_rx =1115;
21911: waveform_sig_rx =1299;
21912: waveform_sig_rx =804;
21913: waveform_sig_rx =1160;
21914: waveform_sig_rx =1300;
21915: waveform_sig_rx =837;
21916: waveform_sig_rx =1190;
21917: waveform_sig_rx =1210;
21918: waveform_sig_rx =1009;
21919: waveform_sig_rx =1041;
21920: waveform_sig_rx =1246;
21921: waveform_sig_rx =1068;
21922: waveform_sig_rx =1047;
21923: waveform_sig_rx =1118;
21924: waveform_sig_rx =1254;
21925: waveform_sig_rx =937;
21926: waveform_sig_rx =1104;
21927: waveform_sig_rx =1298;
21928: waveform_sig_rx =991;
21929: waveform_sig_rx =1040;
21930: waveform_sig_rx =1326;
21931: waveform_sig_rx =1069;
21932: waveform_sig_rx =971;
21933: waveform_sig_rx =1322;
21934: waveform_sig_rx =1117;
21935: waveform_sig_rx =1004;
21936: waveform_sig_rx =1199;
21937: waveform_sig_rx =1235;
21938: waveform_sig_rx =1051;
21939: waveform_sig_rx =1173;
21940: waveform_sig_rx =1085;
21941: waveform_sig_rx =1222;
21942: waveform_sig_rx =1067;
21943: waveform_sig_rx =1211;
21944: waveform_sig_rx =1096;
21945: waveform_sig_rx =1053;
21946: waveform_sig_rx =1372;
21947: waveform_sig_rx =887;
21948: waveform_sig_rx =1256;
21949: waveform_sig_rx =1291;
21950: waveform_sig_rx =871;
21951: waveform_sig_rx =1291;
21952: waveform_sig_rx =1281;
21953: waveform_sig_rx =885;
21954: waveform_sig_rx =1273;
21955: waveform_sig_rx =1275;
21956: waveform_sig_rx =934;
21957: waveform_sig_rx =1239;
21958: waveform_sig_rx =1233;
21959: waveform_sig_rx =1083;
21960: waveform_sig_rx =1074;
21961: waveform_sig_rx =1287;
21962: waveform_sig_rx =1144;
21963: waveform_sig_rx =1042;
21964: waveform_sig_rx =1182;
21965: waveform_sig_rx =1301;
21966: waveform_sig_rx =923;
21967: waveform_sig_rx =1196;
21968: waveform_sig_rx =1296;
21969: waveform_sig_rx =957;
21970: waveform_sig_rx =1144;
21971: waveform_sig_rx =1302;
21972: waveform_sig_rx =1066;
21973: waveform_sig_rx =1048;
21974: waveform_sig_rx =1264;
21975: waveform_sig_rx =1173;
21976: waveform_sig_rx =1030;
21977: waveform_sig_rx =1176;
21978: waveform_sig_rx =1298;
21979: waveform_sig_rx =988;
21980: waveform_sig_rx =1200;
21981: waveform_sig_rx =1112;
21982: waveform_sig_rx =1172;
21983: waveform_sig_rx =1140;
21984: waveform_sig_rx =1237;
21985: waveform_sig_rx =1046;
21986: waveform_sig_rx =1138;
21987: waveform_sig_rx =1335;
21988: waveform_sig_rx =851;
21989: waveform_sig_rx =1303;
21990: waveform_sig_rx =1199;
21991: waveform_sig_rx =897;
21992: waveform_sig_rx =1295;
21993: waveform_sig_rx =1179;
21994: waveform_sig_rx =934;
21995: waveform_sig_rx =1236;
21996: waveform_sig_rx =1213;
21997: waveform_sig_rx =983;
21998: waveform_sig_rx =1146;
21999: waveform_sig_rx =1223;
22000: waveform_sig_rx =1046;
22001: waveform_sig_rx =984;
22002: waveform_sig_rx =1311;
22003: waveform_sig_rx =1054;
22004: waveform_sig_rx =1007;
22005: waveform_sig_rx =1170;
22006: waveform_sig_rx =1216;
22007: waveform_sig_rx =917;
22008: waveform_sig_rx =1173;
22009: waveform_sig_rx =1232;
22010: waveform_sig_rx =940;
22011: waveform_sig_rx =1123;
22012: waveform_sig_rx =1225;
22013: waveform_sig_rx =1044;
22014: waveform_sig_rx =1005;
22015: waveform_sig_rx =1186;
22016: waveform_sig_rx =1178;
22017: waveform_sig_rx =928;
22018: waveform_sig_rx =1155;
22019: waveform_sig_rx =1266;
22020: waveform_sig_rx =853;
22021: waveform_sig_rx =1235;
22022: waveform_sig_rx =1006;
22023: waveform_sig_rx =1101;
22024: waveform_sig_rx =1108;
22025: waveform_sig_rx =1096;
22026: waveform_sig_rx =985;
22027: waveform_sig_rx =1092;
22028: waveform_sig_rx =1165;
22029: waveform_sig_rx =818;
22030: waveform_sig_rx =1215;
22031: waveform_sig_rx =1066;
22032: waveform_sig_rx =878;
22033: waveform_sig_rx =1206;
22034: waveform_sig_rx =1098;
22035: waveform_sig_rx =840;
22036: waveform_sig_rx =1125;
22037: waveform_sig_rx =1135;
22038: waveform_sig_rx =871;
22039: waveform_sig_rx =1047;
22040: waveform_sig_rx =1157;
22041: waveform_sig_rx =915;
22042: waveform_sig_rx =894;
22043: waveform_sig_rx =1251;
22044: waveform_sig_rx =918;
22045: waveform_sig_rx =924;
22046: waveform_sig_rx =1090;
22047: waveform_sig_rx =1073;
22048: waveform_sig_rx =838;
22049: waveform_sig_rx =1057;
22050: waveform_sig_rx =1080;
22051: waveform_sig_rx =872;
22052: waveform_sig_rx =971;
22053: waveform_sig_rx =1126;
22054: waveform_sig_rx =959;
22055: waveform_sig_rx =837;
22056: waveform_sig_rx =1134;
22057: waveform_sig_rx =1017;
22058: waveform_sig_rx =738;
22059: waveform_sig_rx =1105;
22060: waveform_sig_rx =1029;
22061: waveform_sig_rx =742;
22062: waveform_sig_rx =1148;
22063: waveform_sig_rx =783;
22064: waveform_sig_rx =1036;
22065: waveform_sig_rx =931;
22066: waveform_sig_rx =945;
22067: waveform_sig_rx =890;
22068: waveform_sig_rx =896;
22069: waveform_sig_rx =1030;
22070: waveform_sig_rx =695;
22071: waveform_sig_rx =1018;
22072: waveform_sig_rx =963;
22073: waveform_sig_rx =690;
22074: waveform_sig_rx =1049;
22075: waveform_sig_rx =975;
22076: waveform_sig_rx =669;
22077: waveform_sig_rx =987;
22078: waveform_sig_rx =964;
22079: waveform_sig_rx =686;
22080: waveform_sig_rx =890;
22081: waveform_sig_rx =1015;
22082: waveform_sig_rx =695;
22083: waveform_sig_rx =768;
22084: waveform_sig_rx =1069;
22085: waveform_sig_rx =683;
22086: waveform_sig_rx =814;
22087: waveform_sig_rx =883;
22088: waveform_sig_rx =887;
22089: waveform_sig_rx =711;
22090: waveform_sig_rx =836;
22091: waveform_sig_rx =949;
22092: waveform_sig_rx =688;
22093: waveform_sig_rx =739;
22094: waveform_sig_rx =1002;
22095: waveform_sig_rx =698;
22096: waveform_sig_rx =665;
22097: waveform_sig_rx =967;
22098: waveform_sig_rx =724;
22099: waveform_sig_rx =621;
22100: waveform_sig_rx =895;
22101: waveform_sig_rx =797;
22102: waveform_sig_rx =613;
22103: waveform_sig_rx =866;
22104: waveform_sig_rx =613;
22105: waveform_sig_rx =843;
22106: waveform_sig_rx =653;
22107: waveform_sig_rx =780;
22108: waveform_sig_rx =628;
22109: waveform_sig_rx =675;
22110: waveform_sig_rx =836;
22111: waveform_sig_rx =463;
22112: waveform_sig_rx =826;
22113: waveform_sig_rx =731;
22114: waveform_sig_rx =466;
22115: waveform_sig_rx =836;
22116: waveform_sig_rx =760;
22117: waveform_sig_rx =434;
22118: waveform_sig_rx =802;
22119: waveform_sig_rx =752;
22120: waveform_sig_rx =397;
22121: waveform_sig_rx =758;
22122: waveform_sig_rx =752;
22123: waveform_sig_rx =449;
22124: waveform_sig_rx =629;
22125: waveform_sig_rx =719;
22126: waveform_sig_rx =501;
22127: waveform_sig_rx =568;
22128: waveform_sig_rx =589;
22129: waveform_sig_rx =722;
22130: waveform_sig_rx =382;
22131: waveform_sig_rx =639;
22132: waveform_sig_rx =725;
22133: waveform_sig_rx =361;
22134: waveform_sig_rx =583;
22135: waveform_sig_rx =723;
22136: waveform_sig_rx =420;
22137: waveform_sig_rx =469;
22138: waveform_sig_rx =689;
22139: waveform_sig_rx =465;
22140: waveform_sig_rx =396;
22141: waveform_sig_rx =614;
22142: waveform_sig_rx =527;
22143: waveform_sig_rx =364;
22144: waveform_sig_rx =569;
22145: waveform_sig_rx =355;
22146: waveform_sig_rx =591;
22147: waveform_sig_rx =342;
22148: waveform_sig_rx =545;
22149: waveform_sig_rx =332;
22150: waveform_sig_rx =444;
22151: waveform_sig_rx =588;
22152: waveform_sig_rx =172;
22153: waveform_sig_rx =588;
22154: waveform_sig_rx =467;
22155: waveform_sig_rx =153;
22156: waveform_sig_rx =638;
22157: waveform_sig_rx =436;
22158: waveform_sig_rx =143;
22159: waveform_sig_rx =603;
22160: waveform_sig_rx =392;
22161: waveform_sig_rx =179;
22162: waveform_sig_rx =488;
22163: waveform_sig_rx =400;
22164: waveform_sig_rx =230;
22165: waveform_sig_rx =302;
22166: waveform_sig_rx =439;
22167: waveform_sig_rx =293;
22168: waveform_sig_rx =228;
22169: waveform_sig_rx =382;
22170: waveform_sig_rx =419;
22171: waveform_sig_rx =56;
22172: waveform_sig_rx =423;
22173: waveform_sig_rx =373;
22174: waveform_sig_rx =87;
22175: waveform_sig_rx =323;
22176: waveform_sig_rx =384;
22177: waveform_sig_rx =143;
22178: waveform_sig_rx =199;
22179: waveform_sig_rx =384;
22180: waveform_sig_rx =195;
22181: waveform_sig_rx =114;
22182: waveform_sig_rx =309;
22183: waveform_sig_rx =278;
22184: waveform_sig_rx =69;
22185: waveform_sig_rx =258;
22186: waveform_sig_rx =121;
22187: waveform_sig_rx =237;
22188: waveform_sig_rx =85;
22189: waveform_sig_rx =289;
22190: waveform_sig_rx =-31;
22191: waveform_sig_rx =238;
22192: waveform_sig_rx =248;
22193: waveform_sig_rx =-149;
22194: waveform_sig_rx =366;
22195: waveform_sig_rx =80;
22196: waveform_sig_rx =-85;
22197: waveform_sig_rx =337;
22198: waveform_sig_rx =66;
22199: waveform_sig_rx =-75;
22200: waveform_sig_rx =265;
22201: waveform_sig_rx =85;
22202: waveform_sig_rx =-78;
22203: waveform_sig_rx =144;
22204: waveform_sig_rx =135;
22205: waveform_sig_rx =-67;
22206: waveform_sig_rx =-14;
22207: waveform_sig_rx =193;
22208: waveform_sig_rx =-56;
22209: waveform_sig_rx =-95;
22210: waveform_sig_rx =119;
22211: waveform_sig_rx =68;
22212: waveform_sig_rx =-227;
22213: waveform_sig_rx =143;
22214: waveform_sig_rx =21;
22215: waveform_sig_rx =-194;
22216: waveform_sig_rx =21;
22217: waveform_sig_rx =31;
22218: waveform_sig_rx =-133;
22219: waveform_sig_rx =-148;
22220: waveform_sig_rx =55;
22221: waveform_sig_rx =-58;
22222: waveform_sig_rx =-243;
22223: waveform_sig_rx =56;
22224: waveform_sig_rx =-15;
22225: waveform_sig_rx =-295;
22226: waveform_sig_rx =18;
22227: waveform_sig_rx =-210;
22228: waveform_sig_rx =-81;
22229: waveform_sig_rx =-151;
22230: waveform_sig_rx =-67;
22231: waveform_sig_rx =-303;
22232: waveform_sig_rx =3;
22233: waveform_sig_rx =-144;
22234: waveform_sig_rx =-361;
22235: waveform_sig_rx =49;
22236: waveform_sig_rx =-234;
22237: waveform_sig_rx =-338;
22238: waveform_sig_rx =-21;
22239: waveform_sig_rx =-229;
22240: waveform_sig_rx =-391;
22241: waveform_sig_rx =-46;
22242: waveform_sig_rx =-213;
22243: waveform_sig_rx =-375;
22244: waveform_sig_rx =-158;
22245: waveform_sig_rx =-166;
22246: waveform_sig_rx =-381;
22247: waveform_sig_rx =-335;
22248: waveform_sig_rx =-81;
22249: waveform_sig_rx =-391;
22250: waveform_sig_rx =-386;
22251: waveform_sig_rx =-135;
22252: waveform_sig_rx =-313;
22253: waveform_sig_rx =-483;
22254: waveform_sig_rx =-173;
22255: waveform_sig_rx =-318;
22256: waveform_sig_rx =-418;
22257: waveform_sig_rx =-351;
22258: waveform_sig_rx =-215;
22259: waveform_sig_rx =-432;
22260: waveform_sig_rx =-487;
22261: waveform_sig_rx =-151;
22262: waveform_sig_rx =-437;
22263: waveform_sig_rx =-526;
22264: waveform_sig_rx =-202;
22265: waveform_sig_rx =-398;
22266: waveform_sig_rx =-551;
22267: waveform_sig_rx =-301;
22268: waveform_sig_rx =-557;
22269: waveform_sig_rx =-360;
22270: waveform_sig_rx =-474;
22271: waveform_sig_rx =-394;
22272: waveform_sig_rx =-575;
22273: waveform_sig_rx =-329;
22274: waveform_sig_rx =-466;
22275: waveform_sig_rx =-626;
22276: waveform_sig_rx =-287;
22277: waveform_sig_rx =-551;
22278: waveform_sig_rx =-601;
22279: waveform_sig_rx =-334;
22280: waveform_sig_rx =-479;
22281: waveform_sig_rx =-712;
22282: waveform_sig_rx =-371;
22283: waveform_sig_rx =-469;
22284: waveform_sig_rx =-714;
22285: waveform_sig_rx =-433;
22286: waveform_sig_rx =-425;
22287: waveform_sig_rx =-741;
22288: waveform_sig_rx =-560;
22289: waveform_sig_rx =-373;
22290: waveform_sig_rx =-714;
22291: waveform_sig_rx =-608;
22292: waveform_sig_rx =-463;
22293: waveform_sig_rx =-598;
22294: waveform_sig_rx =-705;
22295: waveform_sig_rx =-510;
22296: waveform_sig_rx =-561;
22297: waveform_sig_rx =-724;
22298: waveform_sig_rx =-659;
22299: waveform_sig_rx =-422;
22300: waveform_sig_rx =-780;
22301: waveform_sig_rx =-709;
22302: waveform_sig_rx =-431;
22303: waveform_sig_rx =-778;
22304: waveform_sig_rx =-747;
22305: waveform_sig_rx =-499;
22306: waveform_sig_rx =-700;
22307: waveform_sig_rx =-788;
22308: waveform_sig_rx =-592;
22309: waveform_sig_rx =-824;
22310: waveform_sig_rx =-601;
22311: waveform_sig_rx =-773;
22312: waveform_sig_rx =-655;
22313: waveform_sig_rx =-831;
22314: waveform_sig_rx =-623;
22315: waveform_sig_rx =-731;
22316: waveform_sig_rx =-860;
22317: waveform_sig_rx =-591;
22318: waveform_sig_rx =-741;
22319: waveform_sig_rx =-875;
22320: waveform_sig_rx =-599;
22321: waveform_sig_rx =-688;
22322: waveform_sig_rx =-1031;
22323: waveform_sig_rx =-551;
22324: waveform_sig_rx =-751;
22325: waveform_sig_rx =-1011;
22326: waveform_sig_rx =-604;
22327: waveform_sig_rx =-767;
22328: waveform_sig_rx =-980;
22329: waveform_sig_rx =-785;
22330: waveform_sig_rx =-707;
22331: waveform_sig_rx =-914;
22332: waveform_sig_rx =-899;
22333: waveform_sig_rx =-736;
22334: waveform_sig_rx =-828;
22335: waveform_sig_rx =-1011;
22336: waveform_sig_rx =-715;
22337: waveform_sig_rx =-789;
22338: waveform_sig_rx =-999;
22339: waveform_sig_rx =-861;
22340: waveform_sig_rx =-686;
22341: waveform_sig_rx =-1028;
22342: waveform_sig_rx =-921;
22343: waveform_sig_rx =-641;
22344: waveform_sig_rx =-1018;
22345: waveform_sig_rx =-949;
22346: waveform_sig_rx =-742;
22347: waveform_sig_rx =-921;
22348: waveform_sig_rx =-953;
22349: waveform_sig_rx =-842;
22350: waveform_sig_rx =-1013;
22351: waveform_sig_rx =-808;
22352: waveform_sig_rx =-1028;
22353: waveform_sig_rx =-807;
22354: waveform_sig_rx =-1092;
22355: waveform_sig_rx =-848;
22356: waveform_sig_rx =-899;
22357: waveform_sig_rx =-1148;
22358: waveform_sig_rx =-780;
22359: waveform_sig_rx =-988;
22360: waveform_sig_rx =-1154;
22361: waveform_sig_rx =-725;
22362: waveform_sig_rx =-999;
22363: waveform_sig_rx =-1194;
22364: waveform_sig_rx =-707;
22365: waveform_sig_rx =-1037;
22366: waveform_sig_rx =-1133;
22367: waveform_sig_rx =-823;
22368: waveform_sig_rx =-972;
22369: waveform_sig_rx =-1128;
22370: waveform_sig_rx =-982;
22371: waveform_sig_rx =-874;
22372: waveform_sig_rx =-1080;
22373: waveform_sig_rx =-1080;
22374: waveform_sig_rx =-881;
22375: waveform_sig_rx =-1006;
22376: waveform_sig_rx =-1203;
22377: waveform_sig_rx =-880;
22378: waveform_sig_rx =-985;
22379: waveform_sig_rx =-1205;
22380: waveform_sig_rx =-958;
22381: waveform_sig_rx =-883;
22382: waveform_sig_rx =-1228;
22383: waveform_sig_rx =-1045;
22384: waveform_sig_rx =-895;
22385: waveform_sig_rx =-1158;
22386: waveform_sig_rx =-1125;
22387: waveform_sig_rx =-949;
22388: waveform_sig_rx =-1065;
22389: waveform_sig_rx =-1169;
22390: waveform_sig_rx =-1014;
22391: waveform_sig_rx =-1116;
22392: waveform_sig_rx =-1004;
22393: waveform_sig_rx =-1159;
22394: waveform_sig_rx =-957;
22395: waveform_sig_rx =-1297;
22396: waveform_sig_rx =-903;
22397: waveform_sig_rx =-1087;
22398: waveform_sig_rx =-1278;
22399: waveform_sig_rx =-839;
22400: waveform_sig_rx =-1205;
22401: waveform_sig_rx =-1256;
22402: waveform_sig_rx =-853;
22403: waveform_sig_rx =-1188;
22404: waveform_sig_rx =-1267;
22405: waveform_sig_rx =-861;
22406: waveform_sig_rx =-1199;
22407: waveform_sig_rx =-1230;
22408: waveform_sig_rx =-1008;
22409: waveform_sig_rx =-1085;
22410: waveform_sig_rx =-1256;
22411: waveform_sig_rx =-1117;
22412: waveform_sig_rx =-1001;
22413: waveform_sig_rx =-1208;
22414: waveform_sig_rx =-1217;
22415: waveform_sig_rx =-985;
22416: waveform_sig_rx =-1146;
22417: waveform_sig_rx =-1323;
22418: waveform_sig_rx =-947;
22419: waveform_sig_rx =-1142;
22420: waveform_sig_rx =-1295;
22421: waveform_sig_rx =-1052;
22422: waveform_sig_rx =-1068;
22423: waveform_sig_rx =-1279;
22424: waveform_sig_rx =-1154;
22425: waveform_sig_rx =-1047;
22426: waveform_sig_rx =-1210;
22427: waveform_sig_rx =-1269;
22428: waveform_sig_rx =-990;
22429: waveform_sig_rx =-1154;
22430: waveform_sig_rx =-1262;
22431: waveform_sig_rx =-1057;
22432: waveform_sig_rx =-1217;
22433: waveform_sig_rx =-1090;
22434: waveform_sig_rx =-1195;
22435: waveform_sig_rx =-1058;
22436: waveform_sig_rx =-1347;
22437: waveform_sig_rx =-943;
22438: waveform_sig_rx =-1243;
22439: waveform_sig_rx =-1313;
22440: waveform_sig_rx =-908;
22441: waveform_sig_rx =-1300;
22442: waveform_sig_rx =-1250;
22443: waveform_sig_rx =-940;
22444: waveform_sig_rx =-1290;
22445: waveform_sig_rx =-1259;
22446: waveform_sig_rx =-996;
22447: waveform_sig_rx =-1243;
22448: waveform_sig_rx =-1269;
22449: waveform_sig_rx =-1092;
22450: waveform_sig_rx =-1080;
22451: waveform_sig_rx =-1339;
22452: waveform_sig_rx =-1121;
22453: waveform_sig_rx =-997;
22454: waveform_sig_rx =-1309;
22455: waveform_sig_rx =-1213;
22456: waveform_sig_rx =-1027;
22457: waveform_sig_rx =-1219;
22458: waveform_sig_rx =-1295;
22459: waveform_sig_rx =-1013;
22460: waveform_sig_rx =-1186;
22461: waveform_sig_rx =-1304;
22462: waveform_sig_rx =-1090;
22463: waveform_sig_rx =-1080;
22464: waveform_sig_rx =-1296;
22465: waveform_sig_rx =-1186;
22466: waveform_sig_rx =-1025;
22467: waveform_sig_rx =-1219;
22468: waveform_sig_rx =-1296;
22469: waveform_sig_rx =-962;
22470: waveform_sig_rx =-1202;
22471: waveform_sig_rx =-1269;
22472: waveform_sig_rx =-1016;
22473: waveform_sig_rx =-1271;
22474: waveform_sig_rx =-1049;
22475: waveform_sig_rx =-1165;
22476: waveform_sig_rx =-1099;
22477: waveform_sig_rx =-1302;
22478: waveform_sig_rx =-948;
22479: waveform_sig_rx =-1241;
22480: waveform_sig_rx =-1241;
22481: waveform_sig_rx =-952;
22482: waveform_sig_rx =-1257;
22483: waveform_sig_rx =-1203;
22484: waveform_sig_rx =-961;
22485: waveform_sig_rx =-1204;
22486: waveform_sig_rx =-1271;
22487: waveform_sig_rx =-919;
22488: waveform_sig_rx =-1183;
22489: waveform_sig_rx =-1253;
22490: waveform_sig_rx =-1018;
22491: waveform_sig_rx =-1049;
22492: waveform_sig_rx =-1314;
22493: waveform_sig_rx =-1054;
22494: waveform_sig_rx =-1000;
22495: waveform_sig_rx =-1255;
22496: waveform_sig_rx =-1145;
22497: waveform_sig_rx =-983;
22498: waveform_sig_rx =-1167;
22499: waveform_sig_rx =-1212;
22500: waveform_sig_rx =-942;
22501: waveform_sig_rx =-1129;
22502: waveform_sig_rx =-1189;
22503: waveform_sig_rx =-1050;
22504: waveform_sig_rx =-984;
22505: waveform_sig_rx =-1219;
22506: waveform_sig_rx =-1126;
22507: waveform_sig_rx =-872;
22508: waveform_sig_rx =-1230;
22509: waveform_sig_rx =-1149;
22510: waveform_sig_rx =-839;
22511: waveform_sig_rx =-1221;
22512: waveform_sig_rx =-1081;
22513: waveform_sig_rx =-991;
22514: waveform_sig_rx =-1193;
22515: waveform_sig_rx =-917;
22516: waveform_sig_rx =-1158;
22517: waveform_sig_rx =-981;
22518: waveform_sig_rx =-1197;
22519: waveform_sig_rx =-894;
22520: waveform_sig_rx =-1108;
22521: waveform_sig_rx =-1161;
22522: waveform_sig_rx =-834;
22523: waveform_sig_rx =-1140;
22524: waveform_sig_rx =-1129;
22525: waveform_sig_rx =-793;
22526: waveform_sig_rx =-1127;
22527: waveform_sig_rx =-1140;
22528: waveform_sig_rx =-806;
22529: waveform_sig_rx =-1081;
22530: waveform_sig_rx =-1128;
22531: waveform_sig_rx =-869;
22532: waveform_sig_rx =-945;
22533: waveform_sig_rx =-1222;
22534: waveform_sig_rx =-861;
22535: waveform_sig_rx =-926;
22536: waveform_sig_rx =-1114;
22537: waveform_sig_rx =-977;
22538: waveform_sig_rx =-897;
22539: waveform_sig_rx =-1001;
22540: waveform_sig_rx =-1076;
22541: waveform_sig_rx =-852;
22542: waveform_sig_rx =-934;
22543: waveform_sig_rx =-1114;
22544: waveform_sig_rx =-870;
22545: waveform_sig_rx =-813;
22546: waveform_sig_rx =-1164;
22547: waveform_sig_rx =-896;
22548: waveform_sig_rx =-770;
22549: waveform_sig_rx =-1106;
22550: waveform_sig_rx =-942;
22551: waveform_sig_rx =-756;
22552: waveform_sig_rx =-1018;
22553: waveform_sig_rx =-901;
22554: waveform_sig_rx =-892;
22555: waveform_sig_rx =-953;
22556: waveform_sig_rx =-804;
22557: waveform_sig_rx =-1001;
22558: waveform_sig_rx =-761;
22559: waveform_sig_rx =-1077;
22560: waveform_sig_rx =-686;
22561: waveform_sig_rx =-942;
22562: waveform_sig_rx =-982;
22563: waveform_sig_rx =-651;
22564: waveform_sig_rx =-1007;
22565: waveform_sig_rx =-930;
22566: waveform_sig_rx =-626;
22567: waveform_sig_rx =-962;
22568: waveform_sig_rx =-970;
22569: waveform_sig_rx =-617;
22570: waveform_sig_rx =-905;
22571: waveform_sig_rx =-964;
22572: waveform_sig_rx =-633;
22573: waveform_sig_rx =-824;
22574: waveform_sig_rx =-1008;
22575: waveform_sig_rx =-640;
22576: waveform_sig_rx =-826;
22577: waveform_sig_rx =-841;
22578: waveform_sig_rx =-830;
22579: waveform_sig_rx =-687;
22580: waveform_sig_rx =-741;
22581: waveform_sig_rx =-966;
22582: waveform_sig_rx =-554;
22583: waveform_sig_rx =-770;
22584: waveform_sig_rx =-937;
22585: waveform_sig_rx =-563;
22586: waveform_sig_rx =-728;
22587: waveform_sig_rx =-890;
22588: waveform_sig_rx =-684;
22589: waveform_sig_rx =-612;
22590: waveform_sig_rx =-822;
22591: waveform_sig_rx =-789;
22592: waveform_sig_rx =-527;
22593: waveform_sig_rx =-811;
22594: waveform_sig_rx =-724;
22595: waveform_sig_rx =-673;
22596: waveform_sig_rx =-752;
22597: waveform_sig_rx =-585;
22598: waveform_sig_rx =-755;
22599: waveform_sig_rx =-562;
22600: waveform_sig_rx =-857;
22601: waveform_sig_rx =-453;
22602: waveform_sig_rx =-724;
22603: waveform_sig_rx =-757;
22604: waveform_sig_rx =-387;
22605: waveform_sig_rx =-799;
22606: waveform_sig_rx =-701;
22607: waveform_sig_rx =-337;
22608: waveform_sig_rx =-797;
22609: waveform_sig_rx =-677;
22610: waveform_sig_rx =-359;
22611: waveform_sig_rx =-757;
22612: waveform_sig_rx =-607;
22613: waveform_sig_rx =-457;
22614: waveform_sig_rx =-574;
22615: waveform_sig_rx =-707;
22616: waveform_sig_rx =-483;
22617: waveform_sig_rx =-494;
22618: waveform_sig_rx =-626;
22619: waveform_sig_rx =-604;
22620: waveform_sig_rx =-369;
22621: waveform_sig_rx =-616;
22622: waveform_sig_rx =-662;
22623: waveform_sig_rx =-284;
22624: waveform_sig_rx =-611;
22625: waveform_sig_rx =-630;
22626: waveform_sig_rx =-387;
22627: waveform_sig_rx =-465;
22628: waveform_sig_rx =-612;
22629: waveform_sig_rx =-450;
22630: waveform_sig_rx =-364;
22631: waveform_sig_rx =-589;
22632: waveform_sig_rx =-514;
22633: waveform_sig_rx =-279;
22634: waveform_sig_rx =-552;
22635: waveform_sig_rx =-442;
22636: waveform_sig_rx =-412;
22637: waveform_sig_rx =-456;
22638: waveform_sig_rx =-364;
22639: waveform_sig_rx =-470;
22640: waveform_sig_rx =-317;
22641: waveform_sig_rx =-607;
22642: waveform_sig_rx =-149;
22643: waveform_sig_rx =-522;
22644: waveform_sig_rx =-468;
22645: waveform_sig_rx =-111;
22646: waveform_sig_rx =-592;
22647: waveform_sig_rx =-360;
22648: waveform_sig_rx =-132;
22649: waveform_sig_rx =-555;
22650: waveform_sig_rx =-342;
22651: waveform_sig_rx =-161;
22652: waveform_sig_rx =-441;
22653: waveform_sig_rx =-349;
22654: waveform_sig_rx =-214;
22655: waveform_sig_rx =-250;
22656: waveform_sig_rx =-483;
22657: waveform_sig_rx =-166;
22658: waveform_sig_rx =-188;
22659: waveform_sig_rx =-408;
22660: waveform_sig_rx =-280;
22661: waveform_sig_rx =-93;
22662: waveform_sig_rx =-367;
22663: waveform_sig_rx =-324;
22664: waveform_sig_rx =-61;
22665: waveform_sig_rx =-307;
22666: waveform_sig_rx =-328;
22667: waveform_sig_rx =-100;
22668: waveform_sig_rx =-167;
22669: waveform_sig_rx =-350;
22670: waveform_sig_rx =-135;
22671: waveform_sig_rx =-64;
22672: waveform_sig_rx =-291;
22673: waveform_sig_rx =-226;
22674: waveform_sig_rx =19;
22675: waveform_sig_rx =-258;
22676: waveform_sig_rx =-180;
22677: waveform_sig_rx =-76;
22678: waveform_sig_rx =-185;
22679: waveform_sig_rx =-87;
22680: waveform_sig_rx =-102;
22681: waveform_sig_rx =-101;
22682: waveform_sig_rx =-248;
22683: waveform_sig_rx =135;
22684: waveform_sig_rx =-296;
22685: waveform_sig_rx =-67;
22686: waveform_sig_rx =96;
22687: waveform_sig_rx =-267;
22688: waveform_sig_rx =-49;
22689: waveform_sig_rx =83;
22690: waveform_sig_rx =-182;
22691: waveform_sig_rx =-106;
22692: waveform_sig_rx =164;
22693: waveform_sig_rx =-145;
22694: waveform_sig_rx =-102;
22695: waveform_sig_rx =98;
22696: waveform_sig_rx =3;
22697: waveform_sig_rx =-194;
22698: waveform_sig_rx =136;
22699: waveform_sig_rx =79;
22700: waveform_sig_rx =-136;
22701: waveform_sig_rx =22;
22702: waveform_sig_rx =189;
22703: waveform_sig_rx =-114;
22704: waveform_sig_rx =26;
22705: waveform_sig_rx =205;
22706: waveform_sig_rx =-23;
22707: waveform_sig_rx =-23;
22708: waveform_sig_rx =144;
22709: waveform_sig_rx =178;
22710: waveform_sig_rx =-79;
22711: waveform_sig_rx =158;
22712: waveform_sig_rx =264;
22713: waveform_sig_rx =-80;
22714: waveform_sig_rx =105;
22715: waveform_sig_rx =321;
22716: waveform_sig_rx =-35;
22717: waveform_sig_rx =167;
22718: waveform_sig_rx =158;
22719: waveform_sig_rx =93;
22720: waveform_sig_rx =236;
22721: waveform_sig_rx =142;
22722: waveform_sig_rx =182;
22723: waveform_sig_rx =72;
22724: waveform_sig_rx =382;
22725: waveform_sig_rx =20;
22726: waveform_sig_rx =222;
22727: waveform_sig_rx =334;
22728: waveform_sig_rx =68;
22729: waveform_sig_rx =207;
22730: waveform_sig_rx =386;
22731: waveform_sig_rx =110;
22732: waveform_sig_rx =151;
22733: waveform_sig_rx =478;
22734: waveform_sig_rx =106;
22735: waveform_sig_rx =204;
22736: waveform_sig_rx =437;
22737: waveform_sig_rx =246;
22738: waveform_sig_rx =128;
22739: waveform_sig_rx =473;
22740: waveform_sig_rx =341;
22741: waveform_sig_rx =204;
22742: waveform_sig_rx =329;
22743: waveform_sig_rx =455;
22744: waveform_sig_rx =214;
22745: waveform_sig_rx =295;
22746: waveform_sig_rx =474;
22747: waveform_sig_rx =310;
22748: waveform_sig_rx =240;
22749: waveform_sig_rx =470;
22750: waveform_sig_rx =464;
22751: waveform_sig_rx =157;
22752: waveform_sig_rx =498;
22753: waveform_sig_rx =515;
22754: waveform_sig_rx =194;
22755: waveform_sig_rx =459;
22756: waveform_sig_rx =555;
22757: waveform_sig_rx =269;
22758: waveform_sig_rx =484;
22759: waveform_sig_rx =391;
22760: waveform_sig_rx =418;
22761: waveform_sig_rx =504;
22762: waveform_sig_rx =403;
22763: waveform_sig_rx =516;
22764: waveform_sig_rx =351;
22765: waveform_sig_rx =643;
22766: waveform_sig_rx =342;
22767: waveform_sig_rx =453;
22768: waveform_sig_rx =647;
22769: waveform_sig_rx =346;
22770: waveform_sig_rx =477;
22771: waveform_sig_rx =730;
22772: waveform_sig_rx =348;
22773: waveform_sig_rx =460;
22774: waveform_sig_rx =782;
22775: waveform_sig_rx =324;
22776: waveform_sig_rx =510;
22777: waveform_sig_rx =711;
22778: waveform_sig_rx =476;
22779: waveform_sig_rx =422;
22780: waveform_sig_rx =719;
22781: waveform_sig_rx =575;
22782: waveform_sig_rx =483;
22783: waveform_sig_rx =590;
22784: waveform_sig_rx =739;
22785: waveform_sig_rx =496;
22786: waveform_sig_rx =543;
22787: waveform_sig_rx =774;
22788: waveform_sig_rx =579;
22789: waveform_sig_rx =490;
22790: waveform_sig_rx =796;
22791: waveform_sig_rx =667;
22792: waveform_sig_rx =425;
22793: waveform_sig_rx =818;
22794: waveform_sig_rx =722;
22795: waveform_sig_rx =481;
22796: waveform_sig_rx =736;
22797: waveform_sig_rx =780;
22798: waveform_sig_rx =567;
22799: waveform_sig_rx =728;
22800: waveform_sig_rx =630;
22801: waveform_sig_rx =728;
22802: waveform_sig_rx =688;
22803: waveform_sig_rx =695;
22804: waveform_sig_rx =747;
22805: waveform_sig_rx =556;
22806: waveform_sig_rx =937;
22807: waveform_sig_rx =545;
22808: waveform_sig_rx =705;
22809: waveform_sig_rx =929;
22810: waveform_sig_rx =529;
22811: waveform_sig_rx =769;
22812: waveform_sig_rx =978;
22813: waveform_sig_rx =524;
22814: waveform_sig_rx =774;
22815: waveform_sig_rx =998;
22816: waveform_sig_rx =546;
22817: waveform_sig_rx =804;
22818: waveform_sig_rx =915;
22819: waveform_sig_rx =721;
22820: waveform_sig_rx =674;
22821: waveform_sig_rx =938;
22822: waveform_sig_rx =809;
22823: waveform_sig_rx =718;
22824: waveform_sig_rx =820;
22825: waveform_sig_rx =974;
22826: waveform_sig_rx =696;
22827: waveform_sig_rx =776;
22828: waveform_sig_rx =1014;
22829: waveform_sig_rx =738;
22830: waveform_sig_rx =708;
22831: waveform_sig_rx =1043;
22832: waveform_sig_rx =817;
22833: waveform_sig_rx =693;
22834: waveform_sig_rx =1009;
22835: waveform_sig_rx =897;
22836: waveform_sig_rx =773;
22837: waveform_sig_rx =870;
22838: waveform_sig_rx =1015;
22839: waveform_sig_rx =804;
22840: waveform_sig_rx =880;
22841: waveform_sig_rx =911;
22842: waveform_sig_rx =910;
22843: waveform_sig_rx =870;
22844: waveform_sig_rx =943;
22845: waveform_sig_rx =879;
22846: waveform_sig_rx =821;
22847: waveform_sig_rx =1149;
22848: waveform_sig_rx =694;
22849: waveform_sig_rx =977;
22850: waveform_sig_rx =1076;
22851: waveform_sig_rx =727;
22852: waveform_sig_rx =988;
22853: waveform_sig_rx =1130;
22854: waveform_sig_rx =717;
22855: waveform_sig_rx =985;
22856: waveform_sig_rx =1164;
22857: waveform_sig_rx =731;
22858: waveform_sig_rx =1032;
22859: waveform_sig_rx =1053;
22860: waveform_sig_rx =931;
22861: waveform_sig_rx =874;
22862: waveform_sig_rx =1086;
22863: waveform_sig_rx =1041;
22864: waveform_sig_rx =844;
22865: waveform_sig_rx =1000;
22866: waveform_sig_rx =1198;
22867: waveform_sig_rx =795;
22868: waveform_sig_rx =1036;
22869: waveform_sig_rx =1169;
22870: waveform_sig_rx =873;
22871: waveform_sig_rx =987;
22872: waveform_sig_rx =1130;
22873: waveform_sig_rx =1028;
22874: waveform_sig_rx =892;
22875: waveform_sig_rx =1134;
22876: waveform_sig_rx =1099;
22877: waveform_sig_rx =893;
22878: waveform_sig_rx =1060;
22879: waveform_sig_rx =1213;
22880: waveform_sig_rx =920;
22881: waveform_sig_rx =1085;
22882: waveform_sig_rx =1042;
22883: waveform_sig_rx =1039;
22884: waveform_sig_rx =1071;
22885: waveform_sig_rx =1114;
22886: waveform_sig_rx =1017;
22887: waveform_sig_rx =1000;
22888: waveform_sig_rx =1280;
22889: waveform_sig_rx =816;
22890: waveform_sig_rx =1155;
22891: waveform_sig_rx =1193;
22892: waveform_sig_rx =842;
22893: waveform_sig_rx =1193;
22894: waveform_sig_rx =1206;
22895: waveform_sig_rx =875;
22896: waveform_sig_rx =1140;
22897: waveform_sig_rx =1214;
22898: waveform_sig_rx =921;
22899: waveform_sig_rx =1130;
22900: waveform_sig_rx =1192;
22901: waveform_sig_rx =1096;
22902: waveform_sig_rx =921;
22903: waveform_sig_rx =1273;
22904: waveform_sig_rx =1111;
22905: waveform_sig_rx =931;
22906: waveform_sig_rx =1179;
22907: waveform_sig_rx =1213;
22908: waveform_sig_rx =918;
22909: waveform_sig_rx =1160;
22910: waveform_sig_rx =1198;
22911: waveform_sig_rx =1032;
22912: waveform_sig_rx =1067;
22913: waveform_sig_rx =1232;
22914: waveform_sig_rx =1164;
22915: waveform_sig_rx =953;
22916: waveform_sig_rx =1248;
22917: waveform_sig_rx =1207;
22918: waveform_sig_rx =956;
22919: waveform_sig_rx =1178;
22920: waveform_sig_rx =1294;
22921: waveform_sig_rx =952;
22922: waveform_sig_rx =1198;
22923: waveform_sig_rx =1116;
22924: waveform_sig_rx =1127;
22925: waveform_sig_rx =1135;
22926: waveform_sig_rx =1155;
22927: waveform_sig_rx =1081;
22928: waveform_sig_rx =1108;
22929: waveform_sig_rx =1317;
22930: waveform_sig_rx =893;
22931: waveform_sig_rx =1263;
22932: waveform_sig_rx =1224;
22933: waveform_sig_rx =960;
22934: waveform_sig_rx =1242;
22935: waveform_sig_rx =1258;
22936: waveform_sig_rx =968;
22937: waveform_sig_rx =1149;
22938: waveform_sig_rx =1318;
22939: waveform_sig_rx =973;
22940: waveform_sig_rx =1108;
22941: waveform_sig_rx =1300;
22942: waveform_sig_rx =1056;
22943: waveform_sig_rx =976;
22944: waveform_sig_rx =1346;
22945: waveform_sig_rx =1063;
22946: waveform_sig_rx =1055;
22947: waveform_sig_rx =1209;
22948: waveform_sig_rx =1241;
22949: waveform_sig_rx =994;
22950: waveform_sig_rx =1171;
22951: waveform_sig_rx =1269;
22952: waveform_sig_rx =1036;
22953: waveform_sig_rx =1085;
22954: waveform_sig_rx =1281;
22955: waveform_sig_rx =1149;
22956: waveform_sig_rx =979;
22957: waveform_sig_rx =1273;
22958: waveform_sig_rx =1218;
22959: waveform_sig_rx =929;
22960: waveform_sig_rx =1228;
22961: waveform_sig_rx =1260;
22962: waveform_sig_rx =921;
22963: waveform_sig_rx =1293;
22964: waveform_sig_rx =1027;
22965: waveform_sig_rx =1175;
22966: waveform_sig_rx =1157;
22967: waveform_sig_rx =1127;
22968: waveform_sig_rx =1126;
22969: waveform_sig_rx =1089;
22970: waveform_sig_rx =1298;
22971: waveform_sig_rx =936;
22972: waveform_sig_rx =1213;
22973: waveform_sig_rx =1251;
22974: waveform_sig_rx =929;
22975: waveform_sig_rx =1234;
22976: waveform_sig_rx =1274;
22977: waveform_sig_rx =895;
22978: waveform_sig_rx =1208;
22979: waveform_sig_rx =1272;
22980: waveform_sig_rx =947;
22981: waveform_sig_rx =1142;
22982: waveform_sig_rx =1267;
22983: waveform_sig_rx =1023;
22984: waveform_sig_rx =989;
22985: waveform_sig_rx =1328;
22986: waveform_sig_rx =1030;
22987: waveform_sig_rx =1063;
22988: waveform_sig_rx =1162;
22989: waveform_sig_rx =1197;
22990: waveform_sig_rx =998;
22991: waveform_sig_rx =1106;
22992: waveform_sig_rx =1245;
22993: waveform_sig_rx =1024;
22994: waveform_sig_rx =1009;
22995: waveform_sig_rx =1289;
22996: waveform_sig_rx =1030;
22997: waveform_sig_rx =914;
22998: waveform_sig_rx =1284;
22999: waveform_sig_rx =1080;
23000: waveform_sig_rx =926;
23001: waveform_sig_rx =1189;
23002: waveform_sig_rx =1163;
23003: waveform_sig_rx =927;
23004: waveform_sig_rx =1187;
23005: waveform_sig_rx =952;
23006: waveform_sig_rx =1167;
23007: waveform_sig_rx =1014;
23008: waveform_sig_rx =1088;
23009: waveform_sig_rx =1031;
23010: waveform_sig_rx =978;
23011: waveform_sig_rx =1247;
23012: waveform_sig_rx =819;
23013: waveform_sig_rx =1135;
23014: waveform_sig_rx =1175;
23015: waveform_sig_rx =809;
23016: waveform_sig_rx =1171;
23017: waveform_sig_rx =1147;
23018: waveform_sig_rx =786;
23019: waveform_sig_rx =1131;
23020: waveform_sig_rx =1178;
23021: waveform_sig_rx =832;
23022: waveform_sig_rx =1072;
23023: waveform_sig_rx =1175;
23024: waveform_sig_rx =881;
23025: waveform_sig_rx =948;
23026: waveform_sig_rx =1184;
23027: waveform_sig_rx =916;
23028: waveform_sig_rx =980;
23029: waveform_sig_rx =999;
23030: waveform_sig_rx =1143;
23031: waveform_sig_rx =845;
23032: waveform_sig_rx =986;
23033: waveform_sig_rx =1198;
23034: waveform_sig_rx =796;
23035: waveform_sig_rx =937;
23036: waveform_sig_rx =1168;
23037: waveform_sig_rx =869;
23038: waveform_sig_rx =885;
23039: waveform_sig_rx =1107;
23040: waveform_sig_rx =958;
23041: waveform_sig_rx =842;
23042: waveform_sig_rx =1021;
23043: waveform_sig_rx =1058;
23044: waveform_sig_rx =787;
23045: waveform_sig_rx =1025;
23046: waveform_sig_rx =847;
23047: waveform_sig_rx =993;
23048: waveform_sig_rx =880;
23049: waveform_sig_rx =979;
23050: waveform_sig_rx =858;
23051: waveform_sig_rx =879;
23052: waveform_sig_rx =1099;
23053: waveform_sig_rx =653;
23054: waveform_sig_rx =1026;
23055: waveform_sig_rx =1006;
23056: waveform_sig_rx =630;
23057: waveform_sig_rx =1066;
23058: waveform_sig_rx =988;
23059: waveform_sig_rx =618;
23060: waveform_sig_rx =1040;
23061: waveform_sig_rx =961;
23062: waveform_sig_rx =666;
23063: waveform_sig_rx =976;
23064: waveform_sig_rx =927;
23065: waveform_sig_rx =782;
23066: waveform_sig_rx =780;
23067: waveform_sig_rx =986;
23068: waveform_sig_rx =834;
23069: waveform_sig_rx =729;
23070: waveform_sig_rx =874;
23071: waveform_sig_rx =986;
23072: waveform_sig_rx =585;
23073: waveform_sig_rx =915;
23074: waveform_sig_rx =932;
23075: waveform_sig_rx =622;
23076: waveform_sig_rx =833;
23077: waveform_sig_rx =909;
23078: waveform_sig_rx =734;
23079: waveform_sig_rx =686;
23080: waveform_sig_rx =895;
23081: waveform_sig_rx =789;
23082: waveform_sig_rx =601;
23083: waveform_sig_rx =851;
23084: waveform_sig_rx =860;
23085: waveform_sig_rx =587;
23086: waveform_sig_rx =826;
23087: waveform_sig_rx =648;
23088: waveform_sig_rx =807;
23089: waveform_sig_rx =650;
23090: waveform_sig_rx =814;
23091: waveform_sig_rx =599;
23092: waveform_sig_rx =713;
23093: waveform_sig_rx =890;
23094: waveform_sig_rx =405;
23095: waveform_sig_rx =884;
23096: waveform_sig_rx =737;
23097: waveform_sig_rx =423;
23098: waveform_sig_rx =901;
23099: waveform_sig_rx =667;
23100: waveform_sig_rx =471;
23101: waveform_sig_rx =802;
23102: waveform_sig_rx =693;
23103: waveform_sig_rx =525;
23104: waveform_sig_rx =676;
23105: waveform_sig_rx =735;
23106: waveform_sig_rx =551;
23107: waveform_sig_rx =501;
23108: waveform_sig_rx =812;
23109: waveform_sig_rx =521;
23110: waveform_sig_rx =482;
23111: waveform_sig_rx =695;
23112: waveform_sig_rx =667;
23113: waveform_sig_rx =394;
23114: waveform_sig_rx =673;
23115: waveform_sig_rx =658;
23116: waveform_sig_rx =390;
23117: waveform_sig_rx =570;
23118: waveform_sig_rx =675;
23119: waveform_sig_rx =481;
23120: waveform_sig_rx =440;
23121: waveform_sig_rx =660;
23122: waveform_sig_rx =550;
23123: waveform_sig_rx =351;
23124: waveform_sig_rx =621;
23125: waveform_sig_rx =615;
23126: waveform_sig_rx =301;
23127: waveform_sig_rx =614;
23128: waveform_sig_rx =393;
23129: waveform_sig_rx =523;
23130: waveform_sig_rx =438;
23131: waveform_sig_rx =537;
23132: waveform_sig_rx =320;
23133: waveform_sig_rx =521;
23134: waveform_sig_rx =528;
23135: waveform_sig_rx =187;
23136: waveform_sig_rx =645;
23137: waveform_sig_rx =393;
23138: waveform_sig_rx =258;
23139: waveform_sig_rx =587;
23140: waveform_sig_rx =406;
23141: waveform_sig_rx =256;
23142: waveform_sig_rx =482;
23143: waveform_sig_rx =469;
23144: waveform_sig_rx =217;
23145: waveform_sig_rx =397;
23146: waveform_sig_rx =519;
23147: waveform_sig_rx =213;
23148: waveform_sig_rx =280;
23149: waveform_sig_rx =549;
23150: waveform_sig_rx =243;
23151: waveform_sig_rx =274;
23152: waveform_sig_rx =397;
23153: waveform_sig_rx =377;
23154: waveform_sig_rx =119;
23155: waveform_sig_rx =406;
23156: waveform_sig_rx =366;
23157: waveform_sig_rx =158;
23158: waveform_sig_rx =285;
23159: waveform_sig_rx =397;
23160: waveform_sig_rx =223;
23161: waveform_sig_rx =106;
23162: waveform_sig_rx =408;
23163: waveform_sig_rx =267;
23164: waveform_sig_rx =53;
23165: waveform_sig_rx =399;
23166: waveform_sig_rx =271;
23167: waveform_sig_rx =17;
23168: waveform_sig_rx =376;
23169: waveform_sig_rx =62;
23170: waveform_sig_rx =274;
23171: waveform_sig_rx =159;
23172: waveform_sig_rx =212;
23173: waveform_sig_rx =76;
23174: waveform_sig_rx =218;
23175: waveform_sig_rx =229;
23176: waveform_sig_rx =-61;
23177: waveform_sig_rx =284;
23178: waveform_sig_rx =135;
23179: waveform_sig_rx =-37;
23180: waveform_sig_rx =264;
23181: waveform_sig_rx =159;
23182: waveform_sig_rx =-113;
23183: waveform_sig_rx =231;
23184: waveform_sig_rx =175;
23185: waveform_sig_rx =-129;
23186: waveform_sig_rx =142;
23187: waveform_sig_rx =182;
23188: waveform_sig_rx =-106;
23189: waveform_sig_rx =-5;
23190: waveform_sig_rx =228;
23191: waveform_sig_rx =-72;
23192: waveform_sig_rx =-8;
23193: waveform_sig_rx =108;
23194: waveform_sig_rx =61;
23195: waveform_sig_rx =-153;
23196: waveform_sig_rx =66;
23197: waveform_sig_rx =60;
23198: waveform_sig_rx =-145;
23199: waveform_sig_rx =-73;
23200: waveform_sig_rx =140;
23201: waveform_sig_rx =-140;
23202: waveform_sig_rx =-191;
23203: waveform_sig_rx =155;
23204: waveform_sig_rx =-140;
23205: waveform_sig_rx =-224;
23206: waveform_sig_rx =76;
23207: waveform_sig_rx =-89;
23208: waveform_sig_rx =-226;
23209: waveform_sig_rx =21;
23210: waveform_sig_rx =-242;
23211: waveform_sig_rx =-5;
23212: waveform_sig_rx =-214;
23213: waveform_sig_rx =-65;
23214: waveform_sig_rx =-238;
23215: waveform_sig_rx =-120;
23216: waveform_sig_rx =-69;
23217: waveform_sig_rx =-354;
23218: waveform_sig_rx =-35;
23219: waveform_sig_rx =-141;
23220: waveform_sig_rx =-371;
23221: waveform_sig_rx =-22;
23222: waveform_sig_rx =-137;
23223: waveform_sig_rx =-474;
23224: waveform_sig_rx =-35;
23225: waveform_sig_rx =-178;
23226: waveform_sig_rx =-448;
23227: waveform_sig_rx =-115;
23228: waveform_sig_rx =-173;
23229: waveform_sig_rx =-407;
23230: waveform_sig_rx =-279;
23231: waveform_sig_rx =-112;
23232: waveform_sig_rx =-378;
23233: waveform_sig_rx =-364;
23234: waveform_sig_rx =-221;
23235: waveform_sig_rx =-260;
23236: waveform_sig_rx =-466;
23237: waveform_sig_rx =-235;
23238: waveform_sig_rx =-248;
23239: waveform_sig_rx =-465;
23240: waveform_sig_rx =-381;
23241: waveform_sig_rx =-143;
23242: waveform_sig_rx =-502;
23243: waveform_sig_rx =-449;
23244: waveform_sig_rx =-138;
23245: waveform_sig_rx =-501;
23246: waveform_sig_rx =-441;
23247: waveform_sig_rx =-277;
23248: waveform_sig_rx =-379;
23249: waveform_sig_rx =-480;
23250: waveform_sig_rx =-375;
23251: waveform_sig_rx =-476;
23252: waveform_sig_rx =-331;
23253: waveform_sig_rx =-537;
23254: waveform_sig_rx =-315;
23255: waveform_sig_rx =-586;
23256: waveform_sig_rx =-385;
23257: waveform_sig_rx =-361;
23258: waveform_sig_rx =-700;
23259: waveform_sig_rx =-280;
23260: waveform_sig_rx =-469;
23261: waveform_sig_rx =-687;
23262: waveform_sig_rx =-273;
23263: waveform_sig_rx =-476;
23264: waveform_sig_rx =-733;
23265: waveform_sig_rx =-309;
23266: waveform_sig_rx =-502;
23267: waveform_sig_rx =-718;
23268: waveform_sig_rx =-389;
23269: waveform_sig_rx =-496;
23270: waveform_sig_rx =-697;
23271: waveform_sig_rx =-568;
23272: waveform_sig_rx =-434;
23273: waveform_sig_rx =-642;
23274: waveform_sig_rx =-656;
23275: waveform_sig_rx =-496;
23276: waveform_sig_rx =-525;
23277: waveform_sig_rx =-794;
23278: waveform_sig_rx =-493;
23279: waveform_sig_rx =-520;
23280: waveform_sig_rx =-777;
23281: waveform_sig_rx =-586;
23282: waveform_sig_rx =-453;
23283: waveform_sig_rx =-766;
23284: waveform_sig_rx =-660;
23285: waveform_sig_rx =-470;
23286: waveform_sig_rx =-741;
23287: waveform_sig_rx =-723;
23288: waveform_sig_rx =-588;
23289: waveform_sig_rx =-593;
23290: waveform_sig_rx =-806;
23291: waveform_sig_rx =-628;
23292: waveform_sig_rx =-722;
23293: waveform_sig_rx =-668;
23294: waveform_sig_rx =-751;
23295: waveform_sig_rx =-606;
23296: waveform_sig_rx =-915;
23297: waveform_sig_rx =-572;
23298: waveform_sig_rx =-697;
23299: waveform_sig_rx =-940;
23300: waveform_sig_rx =-527;
23301: waveform_sig_rx =-800;
23302: waveform_sig_rx =-907;
23303: waveform_sig_rx =-550;
23304: waveform_sig_rx =-766;
23305: waveform_sig_rx =-983;
23306: waveform_sig_rx =-569;
23307: waveform_sig_rx =-797;
23308: waveform_sig_rx =-958;
23309: waveform_sig_rx =-651;
23310: waveform_sig_rx =-770;
23311: waveform_sig_rx =-905;
23312: waveform_sig_rx =-836;
23313: waveform_sig_rx =-685;
23314: waveform_sig_rx =-875;
23315: waveform_sig_rx =-949;
23316: waveform_sig_rx =-674;
23317: waveform_sig_rx =-793;
23318: waveform_sig_rx =-1057;
23319: waveform_sig_rx =-639;
23320: waveform_sig_rx =-848;
23321: waveform_sig_rx =-986;
23322: waveform_sig_rx =-787;
23323: waveform_sig_rx =-754;
23324: waveform_sig_rx =-952;
23325: waveform_sig_rx =-945;
23326: waveform_sig_rx =-716;
23327: waveform_sig_rx =-933;
23328: waveform_sig_rx =-1022;
23329: waveform_sig_rx =-736;
23330: waveform_sig_rx =-893;
23331: waveform_sig_rx =-1068;
23332: waveform_sig_rx =-806;
23333: waveform_sig_rx =-1015;
23334: waveform_sig_rx =-870;
23335: waveform_sig_rx =-981;
23336: waveform_sig_rx =-850;
23337: waveform_sig_rx =-1095;
23338: waveform_sig_rx =-801;
23339: waveform_sig_rx =-942;
23340: waveform_sig_rx =-1121;
23341: waveform_sig_rx =-713;
23342: waveform_sig_rx =-1023;
23343: waveform_sig_rx =-1106;
23344: waveform_sig_rx =-742;
23345: waveform_sig_rx =-1027;
23346: waveform_sig_rx =-1133;
23347: waveform_sig_rx =-783;
23348: waveform_sig_rx =-1026;
23349: waveform_sig_rx =-1110;
23350: waveform_sig_rx =-926;
23351: waveform_sig_rx =-899;
23352: waveform_sig_rx =-1116;
23353: waveform_sig_rx =-1055;
23354: waveform_sig_rx =-799;
23355: waveform_sig_rx =-1164;
23356: waveform_sig_rx =-1085;
23357: waveform_sig_rx =-841;
23358: waveform_sig_rx =-1091;
23359: waveform_sig_rx =-1141;
23360: waveform_sig_rx =-897;
23361: waveform_sig_rx =-1024;
23362: waveform_sig_rx =-1127;
23363: waveform_sig_rx =-1043;
23364: waveform_sig_rx =-873;
23365: waveform_sig_rx =-1175;
23366: waveform_sig_rx =-1133;
23367: waveform_sig_rx =-846;
23368: waveform_sig_rx =-1156;
23369: waveform_sig_rx =-1169;
23370: waveform_sig_rx =-896;
23371: waveform_sig_rx =-1077;
23372: waveform_sig_rx =-1188;
23373: waveform_sig_rx =-968;
23374: waveform_sig_rx =-1186;
23375: waveform_sig_rx =-1017;
23376: waveform_sig_rx =-1120;
23377: waveform_sig_rx =-1012;
23378: waveform_sig_rx =-1228;
23379: waveform_sig_rx =-924;
23380: waveform_sig_rx =-1143;
23381: waveform_sig_rx =-1243;
23382: waveform_sig_rx =-911;
23383: waveform_sig_rx =-1215;
23384: waveform_sig_rx =-1184;
23385: waveform_sig_rx =-953;
23386: waveform_sig_rx =-1129;
23387: waveform_sig_rx =-1278;
23388: waveform_sig_rx =-950;
23389: waveform_sig_rx =-1101;
23390: waveform_sig_rx =-1283;
23391: waveform_sig_rx =-1011;
23392: waveform_sig_rx =-1009;
23393: waveform_sig_rx =-1316;
23394: waveform_sig_rx =-1059;
23395: waveform_sig_rx =-963;
23396: waveform_sig_rx =-1277;
23397: waveform_sig_rx =-1145;
23398: waveform_sig_rx =-1048;
23399: waveform_sig_rx =-1145;
23400: waveform_sig_rx =-1255;
23401: waveform_sig_rx =-1023;
23402: waveform_sig_rx =-1092;
23403: waveform_sig_rx =-1280;
23404: waveform_sig_rx =-1125;
23405: waveform_sig_rx =-1004;
23406: waveform_sig_rx =-1280;
23407: waveform_sig_rx =-1186;
23408: waveform_sig_rx =-953;
23409: waveform_sig_rx =-1260;
23410: waveform_sig_rx =-1264;
23411: waveform_sig_rx =-955;
23412: waveform_sig_rx =-1191;
23413: waveform_sig_rx =-1268;
23414: waveform_sig_rx =-1030;
23415: waveform_sig_rx =-1286;
23416: waveform_sig_rx =-1040;
23417: waveform_sig_rx =-1234;
23418: waveform_sig_rx =-1094;
23419: waveform_sig_rx =-1292;
23420: waveform_sig_rx =-1036;
23421: waveform_sig_rx =-1167;
23422: waveform_sig_rx =-1273;
23423: waveform_sig_rx =-994;
23424: waveform_sig_rx =-1195;
23425: waveform_sig_rx =-1292;
23426: waveform_sig_rx =-973;
23427: waveform_sig_rx =-1178;
23428: waveform_sig_rx =-1395;
23429: waveform_sig_rx =-910;
23430: waveform_sig_rx =-1207;
23431: waveform_sig_rx =-1329;
23432: waveform_sig_rx =-985;
23433: waveform_sig_rx =-1138;
23434: waveform_sig_rx =-1328;
23435: waveform_sig_rx =-1112;
23436: waveform_sig_rx =-1063;
23437: waveform_sig_rx =-1271;
23438: waveform_sig_rx =-1193;
23439: waveform_sig_rx =-1060;
23440: waveform_sig_rx =-1168;
23441: waveform_sig_rx =-1289;
23442: waveform_sig_rx =-1046;
23443: waveform_sig_rx =-1100;
23444: waveform_sig_rx =-1293;
23445: waveform_sig_rx =-1130;
23446: waveform_sig_rx =-990;
23447: waveform_sig_rx =-1352;
23448: waveform_sig_rx =-1174;
23449: waveform_sig_rx =-950;
23450: waveform_sig_rx =-1311;
23451: waveform_sig_rx =-1186;
23452: waveform_sig_rx =-996;
23453: waveform_sig_rx =-1215;
23454: waveform_sig_rx =-1166;
23455: waveform_sig_rx =-1114;
23456: waveform_sig_rx =-1220;
23457: waveform_sig_rx =-1021;
23458: waveform_sig_rx =-1261;
23459: waveform_sig_rx =-1010;
23460: waveform_sig_rx =-1304;
23461: waveform_sig_rx =-1012;
23462: waveform_sig_rx =-1123;
23463: waveform_sig_rx =-1302;
23464: waveform_sig_rx =-917;
23465: waveform_sig_rx =-1216;
23466: waveform_sig_rx =-1289;
23467: waveform_sig_rx =-878;
23468: waveform_sig_rx =-1226;
23469: waveform_sig_rx =-1307;
23470: waveform_sig_rx =-889;
23471: waveform_sig_rx =-1209;
23472: waveform_sig_rx =-1253;
23473: waveform_sig_rx =-952;
23474: waveform_sig_rx =-1093;
23475: waveform_sig_rx =-1302;
23476: waveform_sig_rx =-1000;
23477: waveform_sig_rx =-1052;
23478: waveform_sig_rx =-1197;
23479: waveform_sig_rx =-1143;
23480: waveform_sig_rx =-1046;
23481: waveform_sig_rx =-1062;
23482: waveform_sig_rx =-1296;
23483: waveform_sig_rx =-949;
23484: waveform_sig_rx =-1054;
23485: waveform_sig_rx =-1320;
23486: waveform_sig_rx =-971;
23487: waveform_sig_rx =-978;
23488: waveform_sig_rx =-1278;
23489: waveform_sig_rx =-1025;
23490: waveform_sig_rx =-952;
23491: waveform_sig_rx =-1187;
23492: waveform_sig_rx =-1126;
23493: waveform_sig_rx =-943;
23494: waveform_sig_rx =-1104;
23495: waveform_sig_rx =-1109;
23496: waveform_sig_rx =-1031;
23497: waveform_sig_rx =-1118;
23498: waveform_sig_rx =-974;
23499: waveform_sig_rx =-1151;
23500: waveform_sig_rx =-893;
23501: waveform_sig_rx =-1261;
23502: waveform_sig_rx =-868;
23503: waveform_sig_rx =-1067;
23504: waveform_sig_rx =-1244;
23505: waveform_sig_rx =-778;
23506: waveform_sig_rx =-1166;
23507: waveform_sig_rx =-1154;
23508: waveform_sig_rx =-765;
23509: waveform_sig_rx =-1171;
23510: waveform_sig_rx =-1129;
23511: waveform_sig_rx =-761;
23512: waveform_sig_rx =-1136;
23513: waveform_sig_rx =-1093;
23514: waveform_sig_rx =-872;
23515: waveform_sig_rx =-973;
23516: waveform_sig_rx =-1141;
23517: waveform_sig_rx =-934;
23518: waveform_sig_rx =-898;
23519: waveform_sig_rx =-1033;
23520: waveform_sig_rx =-1054;
23521: waveform_sig_rx =-827;
23522: waveform_sig_rx =-968;
23523: waveform_sig_rx =-1166;
23524: waveform_sig_rx =-729;
23525: waveform_sig_rx =-983;
23526: waveform_sig_rx =-1122;
23527: waveform_sig_rx =-798;
23528: waveform_sig_rx =-918;
23529: waveform_sig_rx =-1059;
23530: waveform_sig_rx =-923;
23531: waveform_sig_rx =-808;
23532: waveform_sig_rx =-998;
23533: waveform_sig_rx =-1007;
23534: waveform_sig_rx =-727;
23535: waveform_sig_rx =-963;
23536: waveform_sig_rx =-969;
23537: waveform_sig_rx =-851;
23538: waveform_sig_rx =-945;
23539: waveform_sig_rx =-824;
23540: waveform_sig_rx =-949;
23541: waveform_sig_rx =-761;
23542: waveform_sig_rx =-1102;
23543: waveform_sig_rx =-639;
23544: waveform_sig_rx =-961;
23545: waveform_sig_rx =-1018;
23546: waveform_sig_rx =-563;
23547: waveform_sig_rx =-1061;
23548: waveform_sig_rx =-893;
23549: waveform_sig_rx =-590;
23550: waveform_sig_rx =-1026;
23551: waveform_sig_rx =-874;
23552: waveform_sig_rx =-662;
23553: waveform_sig_rx =-918;
23554: waveform_sig_rx =-887;
23555: waveform_sig_rx =-741;
23556: waveform_sig_rx =-727;
23557: waveform_sig_rx =-1002;
23558: waveform_sig_rx =-730;
23559: waveform_sig_rx =-690;
23560: waveform_sig_rx =-922;
23561: waveform_sig_rx =-825;
23562: waveform_sig_rx =-647;
23563: waveform_sig_rx =-826;
23564: waveform_sig_rx =-907;
23565: waveform_sig_rx =-572;
23566: waveform_sig_rx =-821;
23567: waveform_sig_rx =-882;
23568: waveform_sig_rx =-623;
23569: waveform_sig_rx =-685;
23570: waveform_sig_rx =-836;
23571: waveform_sig_rx =-741;
23572: waveform_sig_rx =-601;
23573: waveform_sig_rx =-797;
23574: waveform_sig_rx =-832;
23575: waveform_sig_rx =-495;
23576: waveform_sig_rx =-795;
23577: waveform_sig_rx =-771;
23578: waveform_sig_rx =-592;
23579: waveform_sig_rx =-792;
23580: waveform_sig_rx =-601;
23581: waveform_sig_rx =-701;
23582: waveform_sig_rx =-613;
23583: waveform_sig_rx =-823;
23584: waveform_sig_rx =-425;
23585: waveform_sig_rx =-797;
23586: waveform_sig_rx =-695;
23587: waveform_sig_rx =-437;
23588: waveform_sig_rx =-815;
23589: waveform_sig_rx =-627;
23590: waveform_sig_rx =-453;
23591: waveform_sig_rx =-725;
23592: waveform_sig_rx =-668;
23593: waveform_sig_rx =-432;
23594: waveform_sig_rx =-629;
23595: waveform_sig_rx =-672;
23596: waveform_sig_rx =-467;
23597: waveform_sig_rx =-507;
23598: waveform_sig_rx =-772;
23599: waveform_sig_rx =-432;
23600: waveform_sig_rx =-472;
23601: waveform_sig_rx =-692;
23602: waveform_sig_rx =-533;
23603: waveform_sig_rx =-388;
23604: waveform_sig_rx =-606;
23605: waveform_sig_rx =-613;
23606: waveform_sig_rx =-358;
23607: waveform_sig_rx =-558;
23608: waveform_sig_rx =-610;
23609: waveform_sig_rx =-421;
23610: waveform_sig_rx =-393;
23611: waveform_sig_rx =-615;
23612: waveform_sig_rx =-492;
23613: waveform_sig_rx =-278;
23614: waveform_sig_rx =-630;
23615: waveform_sig_rx =-535;
23616: waveform_sig_rx =-215;
23617: waveform_sig_rx =-602;
23618: waveform_sig_rx =-439;
23619: waveform_sig_rx =-355;
23620: waveform_sig_rx =-514;
23621: waveform_sig_rx =-291;
23622: waveform_sig_rx =-474;
23623: waveform_sig_rx =-346;
23624: waveform_sig_rx =-524;
23625: waveform_sig_rx =-200;
23626: waveform_sig_rx =-501;
23627: waveform_sig_rx =-424;
23628: waveform_sig_rx =-214;
23629: waveform_sig_rx =-508;
23630: waveform_sig_rx =-402;
23631: waveform_sig_rx =-166;
23632: waveform_sig_rx =-448;
23633: waveform_sig_rx =-448;
23634: waveform_sig_rx =-110;
23635: waveform_sig_rx =-394;
23636: waveform_sig_rx =-431;
23637: waveform_sig_rx =-160;
23638: waveform_sig_rx =-276;
23639: waveform_sig_rx =-518;
23640: waveform_sig_rx =-124;
23641: waveform_sig_rx =-235;
23642: waveform_sig_rx =-403;
23643: waveform_sig_rx =-255;
23644: waveform_sig_rx =-176;
23645: waveform_sig_rx =-316;
23646: waveform_sig_rx =-343;
23647: waveform_sig_rx =-112;
23648: waveform_sig_rx =-232;
23649: waveform_sig_rx =-358;
23650: waveform_sig_rx =-129;
23651: waveform_sig_rx =-88;
23652: waveform_sig_rx =-408;
23653: waveform_sig_rx =-136;
23654: waveform_sig_rx =-17;
23655: waveform_sig_rx =-378;
23656: waveform_sig_rx =-159;
23657: waveform_sig_rx =5;
23658: waveform_sig_rx =-280;
23659: waveform_sig_rx =-125;
23660: waveform_sig_rx =-158;
23661: waveform_sig_rx =-191;
23662: waveform_sig_rx =-56;
23663: waveform_sig_rx =-210;
23664: waveform_sig_rx =-40;
23665: waveform_sig_rx =-266;
23666: waveform_sig_rx =75;
23667: waveform_sig_rx =-200;
23668: waveform_sig_rx =-168;
23669: waveform_sig_rx =99;
23670: waveform_sig_rx =-206;
23671: waveform_sig_rx =-129;
23672: waveform_sig_rx =169;
23673: waveform_sig_rx =-190;
23674: waveform_sig_rx =-162;
23675: waveform_sig_rx =224;
23676: waveform_sig_rx =-172;
23677: waveform_sig_rx =-101;
23678: waveform_sig_rx =185;
23679: waveform_sig_rx =-31;
23680: waveform_sig_rx =-160;
23681: waveform_sig_rx =165;
23682: waveform_sig_rx =28;
23683: waveform_sig_rx =-36;
23684: waveform_sig_rx =12;
23685: waveform_sig_rx =174;
23686: waveform_sig_rx =-3;
23687: waveform_sig_rx =-75;
23688: waveform_sig_rx =252;
23689: waveform_sig_rx =35;
23690: waveform_sig_rx =-84;
23691: waveform_sig_rx =218;
23692: waveform_sig_rx =165;
23693: waveform_sig_rx =-128;
23694: waveform_sig_rx =217;
23695: waveform_sig_rx =213;
23696: waveform_sig_rx =-49;
23697: waveform_sig_rx =151;
23698: waveform_sig_rx =258;
23699: waveform_sig_rx =37;
23700: waveform_sig_rx =159;
23701: waveform_sig_rx =125;
23702: waveform_sig_rx =167;
23703: waveform_sig_rx =190;
23704: waveform_sig_rx =127;
23705: waveform_sig_rx =268;
23706: waveform_sig_rx =-9;
23707: waveform_sig_rx =421;
23708: waveform_sig_rx =73;
23709: waveform_sig_rx =113;
23710: waveform_sig_rx =448;
23711: waveform_sig_rx =28;
23712: waveform_sig_rx =188;
23713: waveform_sig_rx =479;
23714: waveform_sig_rx =36;
23715: waveform_sig_rx =193;
23716: waveform_sig_rx =493;
23717: waveform_sig_rx =69;
23718: waveform_sig_rx =243;
23719: waveform_sig_rx =422;
23720: waveform_sig_rx =230;
23721: waveform_sig_rx =149;
23722: waveform_sig_rx =404;
23723: waveform_sig_rx =327;
23724: waveform_sig_rx =223;
23725: waveform_sig_rx =264;
23726: waveform_sig_rx =505;
23727: waveform_sig_rx =236;
23728: waveform_sig_rx =205;
23729: waveform_sig_rx =567;
23730: waveform_sig_rx =293;
23731: waveform_sig_rx =220;
23732: waveform_sig_rx =553;
23733: waveform_sig_rx =385;
23734: waveform_sig_rx =217;
23735: waveform_sig_rx =493;
23736: waveform_sig_rx =443;
23737: waveform_sig_rx =297;
23738: waveform_sig_rx =378;
23739: waveform_sig_rx =552;
23740: waveform_sig_rx =352;
23741: waveform_sig_rx =375;
23742: waveform_sig_rx =465;
23743: waveform_sig_rx =443;
23744: waveform_sig_rx =435;
23745: waveform_sig_rx =484;
23746: waveform_sig_rx =485;
23747: waveform_sig_rx =308;
23748: waveform_sig_rx =738;
23749: waveform_sig_rx =270;
23750: waveform_sig_rx =479;
23751: waveform_sig_rx =695;
23752: waveform_sig_rx =284;
23753: waveform_sig_rx =513;
23754: waveform_sig_rx =714;
23755: waveform_sig_rx =312;
23756: waveform_sig_rx =495;
23757: waveform_sig_rx =749;
23758: waveform_sig_rx =339;
23759: waveform_sig_rx =555;
23760: waveform_sig_rx =644;
23761: waveform_sig_rx =525;
23762: waveform_sig_rx =431;
23763: waveform_sig_rx =641;
23764: waveform_sig_rx =654;
23765: waveform_sig_rx =440;
23766: waveform_sig_rx =551;
23767: waveform_sig_rx =808;
23768: waveform_sig_rx =416;
23769: waveform_sig_rx =565;
23770: waveform_sig_rx =807;
23771: waveform_sig_rx =467;
23772: waveform_sig_rx =564;
23773: waveform_sig_rx =747;
23774: waveform_sig_rx =654;
23775: waveform_sig_rx =510;
23776: waveform_sig_rx =719;
23777: waveform_sig_rx =755;
23778: waveform_sig_rx =542;
23779: waveform_sig_rx =627;
23780: waveform_sig_rx =866;
23781: waveform_sig_rx =563;
23782: waveform_sig_rx =657;
23783: waveform_sig_rx =750;
23784: waveform_sig_rx =652;
23785: waveform_sig_rx =734;
23786: waveform_sig_rx =752;
23787: waveform_sig_rx =692;
23788: waveform_sig_rx =612;
23789: waveform_sig_rx =945;
23790: waveform_sig_rx =510;
23791: waveform_sig_rx =782;
23792: waveform_sig_rx =891;
23793: waveform_sig_rx =538;
23794: waveform_sig_rx =804;
23795: waveform_sig_rx =934;
23796: waveform_sig_rx =553;
23797: waveform_sig_rx =784;
23798: waveform_sig_rx =948;
23799: waveform_sig_rx =615;
23800: waveform_sig_rx =794;
23801: waveform_sig_rx =854;
23802: waveform_sig_rx =834;
23803: waveform_sig_rx =605;
23804: waveform_sig_rx =945;
23805: waveform_sig_rx =899;
23806: waveform_sig_rx =613;
23807: waveform_sig_rx =886;
23808: waveform_sig_rx =959;
23809: waveform_sig_rx =650;
23810: waveform_sig_rx =882;
23811: waveform_sig_rx =914;
23812: waveform_sig_rx =781;
23813: waveform_sig_rx =768;
23814: waveform_sig_rx =958;
23815: waveform_sig_rx =941;
23816: waveform_sig_rx =663;
23817: waveform_sig_rx =991;
23818: waveform_sig_rx =964;
23819: waveform_sig_rx =693;
23820: waveform_sig_rx =920;
23821: waveform_sig_rx =1041;
23822: waveform_sig_rx =754;
23823: waveform_sig_rx =906;
23824: waveform_sig_rx =923;
23825: waveform_sig_rx =865;
23826: waveform_sig_rx =923;
23827: waveform_sig_rx =939;
23828: waveform_sig_rx =862;
23829: waveform_sig_rx =853;
23830: waveform_sig_rx =1119;
23831: waveform_sig_rx =691;
23832: waveform_sig_rx =1026;
23833: waveform_sig_rx =1031;
23834: waveform_sig_rx =769;
23835: waveform_sig_rx =1005;
23836: waveform_sig_rx =1082;
23837: waveform_sig_rx =828;
23838: waveform_sig_rx =891;
23839: waveform_sig_rx =1170;
23840: waveform_sig_rx =816;
23841: waveform_sig_rx =905;
23842: waveform_sig_rx =1154;
23843: waveform_sig_rx =926;
23844: waveform_sig_rx =783;
23845: waveform_sig_rx =1184;
23846: waveform_sig_rx =958;
23847: waveform_sig_rx =872;
23848: waveform_sig_rx =1053;
23849: waveform_sig_rx =1083;
23850: waveform_sig_rx =883;
23851: waveform_sig_rx =982;
23852: waveform_sig_rx =1135;
23853: waveform_sig_rx =951;
23854: waveform_sig_rx =869;
23855: waveform_sig_rx =1153;
23856: waveform_sig_rx =1069;
23857: waveform_sig_rx =813;
23858: waveform_sig_rx =1157;
23859: waveform_sig_rx =1119;
23860: waveform_sig_rx =850;
23861: waveform_sig_rx =1059;
23862: waveform_sig_rx =1186;
23863: waveform_sig_rx =848;
23864: waveform_sig_rx =1107;
23865: waveform_sig_rx =1020;
23866: waveform_sig_rx =1022;
23867: waveform_sig_rx =1115;
23868: waveform_sig_rx =1034;
23869: waveform_sig_rx =1045;
23870: waveform_sig_rx =999;
23871: waveform_sig_rx =1211;
23872: waveform_sig_rx =892;
23873: waveform_sig_rx =1108;
23874: waveform_sig_rx =1194;
23875: waveform_sig_rx =945;
23876: waveform_sig_rx =1075;
23877: waveform_sig_rx =1298;
23878: waveform_sig_rx =892;
23879: waveform_sig_rx =1058;
23880: waveform_sig_rx =1345;
23881: waveform_sig_rx =864;
23882: waveform_sig_rx =1113;
23883: waveform_sig_rx =1270;
23884: waveform_sig_rx =997;
23885: waveform_sig_rx =986;
23886: waveform_sig_rx =1270;
23887: waveform_sig_rx =1076;
23888: waveform_sig_rx =1038;
23889: waveform_sig_rx =1122;
23890: waveform_sig_rx =1228;
23891: waveform_sig_rx =975;
23892: waveform_sig_rx =1096;
23893: waveform_sig_rx =1274;
23894: waveform_sig_rx =1039;
23895: waveform_sig_rx =1003;
23896: waveform_sig_rx =1278;
23897: waveform_sig_rx =1138;
23898: waveform_sig_rx =896;
23899: waveform_sig_rx =1287;
23900: waveform_sig_rx =1169;
23901: waveform_sig_rx =931;
23902: waveform_sig_rx =1224;
23903: waveform_sig_rx =1215;
23904: waveform_sig_rx =972;
23905: waveform_sig_rx =1221;
23906: waveform_sig_rx =1029;
23907: waveform_sig_rx =1205;
23908: waveform_sig_rx =1120;
23909: waveform_sig_rx =1101;
23910: waveform_sig_rx =1182;
23911: waveform_sig_rx =1007;
23912: waveform_sig_rx =1370;
23913: waveform_sig_rx =965;
23914: waveform_sig_rx =1146;
23915: waveform_sig_rx =1340;
23916: waveform_sig_rx =896;
23917: waveform_sig_rx =1200;
23918: waveform_sig_rx =1334;
23919: waveform_sig_rx =879;
23920: waveform_sig_rx =1206;
23921: waveform_sig_rx =1328;
23922: waveform_sig_rx =938;
23923: waveform_sig_rx =1183;
23924: waveform_sig_rx =1273;
23925: waveform_sig_rx =1066;
23926: waveform_sig_rx =1035;
23927: waveform_sig_rx =1328;
23928: waveform_sig_rx =1112;
23929: waveform_sig_rx =1057;
23930: waveform_sig_rx =1132;
23931: waveform_sig_rx =1268;
23932: waveform_sig_rx =1005;
23933: waveform_sig_rx =1096;
23934: waveform_sig_rx =1339;
23935: waveform_sig_rx =1027;
23936: waveform_sig_rx =1028;
23937: waveform_sig_rx =1363;
23938: waveform_sig_rx =1074;
23939: waveform_sig_rx =1013;
23940: waveform_sig_rx =1320;
23941: waveform_sig_rx =1137;
23942: waveform_sig_rx =1060;
23943: waveform_sig_rx =1168;
23944: waveform_sig_rx =1267;
23945: waveform_sig_rx =1031;
23946: waveform_sig_rx =1167;
23947: waveform_sig_rx =1105;
23948: waveform_sig_rx =1183;
23949: waveform_sig_rx =1089;
23950: waveform_sig_rx =1189;
23951: waveform_sig_rx =1102;
23952: waveform_sig_rx =1027;
23953: waveform_sig_rx =1377;
23954: waveform_sig_rx =865;
23955: waveform_sig_rx =1216;
23956: waveform_sig_rx =1279;
23957: waveform_sig_rx =858;
23958: waveform_sig_rx =1256;
23959: waveform_sig_rx =1251;
23960: waveform_sig_rx =849;
23961: waveform_sig_rx =1223;
23962: waveform_sig_rx =1258;
23963: waveform_sig_rx =927;
23964: waveform_sig_rx =1172;
23965: waveform_sig_rx =1212;
23966: waveform_sig_rx =1059;
23967: waveform_sig_rx =990;
23968: waveform_sig_rx =1269;
23969: waveform_sig_rx =1094;
23970: waveform_sig_rx =1027;
23971: waveform_sig_rx =1124;
23972: waveform_sig_rx =1279;
23973: waveform_sig_rx =914;
23974: waveform_sig_rx =1127;
23975: waveform_sig_rx =1285;
23976: waveform_sig_rx =915;
23977: waveform_sig_rx =1084;
23978: waveform_sig_rx =1262;
23979: waveform_sig_rx =1030;
23980: waveform_sig_rx =1009;
23981: waveform_sig_rx =1198;
23982: waveform_sig_rx =1116;
23983: waveform_sig_rx =973;
23984: waveform_sig_rx =1089;
23985: waveform_sig_rx =1245;
23986: waveform_sig_rx =913;
23987: waveform_sig_rx =1130;
23988: waveform_sig_rx =1057;
23989: waveform_sig_rx =1072;
23990: waveform_sig_rx =1058;
23991: waveform_sig_rx =1131;
23992: waveform_sig_rx =968;
23993: waveform_sig_rx =1024;
23994: waveform_sig_rx =1272;
23995: waveform_sig_rx =767;
23996: waveform_sig_rx =1205;
23997: waveform_sig_rx =1134;
23998: waveform_sig_rx =797;
23999: waveform_sig_rx =1196;
24000: waveform_sig_rx =1115;
24001: waveform_sig_rx =836;
24002: waveform_sig_rx =1140;
24003: waveform_sig_rx =1139;
24004: waveform_sig_rx =890;
24005: waveform_sig_rx =1059;
24006: waveform_sig_rx =1113;
24007: waveform_sig_rx =990;
24008: waveform_sig_rx =867;
24009: waveform_sig_rx =1190;
24010: waveform_sig_rx =978;
24011: waveform_sig_rx =876;
24012: waveform_sig_rx =1070;
24013: waveform_sig_rx =1105;
24014: waveform_sig_rx =780;
24015: waveform_sig_rx =1061;
24016: waveform_sig_rx =1104;
24017: waveform_sig_rx =824;
24018: waveform_sig_rx =1006;
24019: waveform_sig_rx =1086;
24020: waveform_sig_rx =945;
24021: waveform_sig_rx =852;
24022: waveform_sig_rx =1059;
24023: waveform_sig_rx =1054;
24024: waveform_sig_rx =763;
24025: waveform_sig_rx =1031;
24026: waveform_sig_rx =1126;
24027: waveform_sig_rx =725;
24028: waveform_sig_rx =1093;
24029: waveform_sig_rx =864;
24030: waveform_sig_rx =953;
24031: waveform_sig_rx =951;
24032: waveform_sig_rx =960;
24033: waveform_sig_rx =844;
24034: waveform_sig_rx =922;
24035: waveform_sig_rx =1072;
24036: waveform_sig_rx =670;
24037: waveform_sig_rx =1063;
24038: waveform_sig_rx =928;
24039: waveform_sig_rx =683;
24040: waveform_sig_rx =1027;
24041: waveform_sig_rx =932;
24042: waveform_sig_rx =704;
24043: waveform_sig_rx =925;
24044: waveform_sig_rx =980;
24045: waveform_sig_rx =725;
24046: waveform_sig_rx =835;
24047: waveform_sig_rx =1008;
24048: waveform_sig_rx =753;
24049: waveform_sig_rx =694;
24050: waveform_sig_rx =1063;
24051: waveform_sig_rx =740;
24052: waveform_sig_rx =726;
24053: waveform_sig_rx =898;
24054: waveform_sig_rx =893;
24055: waveform_sig_rx =634;
24056: waveform_sig_rx =879;
24057: waveform_sig_rx =891;
24058: waveform_sig_rx =686;
24059: waveform_sig_rx =777;
24060: waveform_sig_rx =892;
24061: waveform_sig_rx =792;
24062: waveform_sig_rx =602;
24063: waveform_sig_rx =920;
24064: waveform_sig_rx =818;
24065: waveform_sig_rx =513;
24066: waveform_sig_rx =911;
24067: waveform_sig_rx =836;
24068: waveform_sig_rx =540;
24069: waveform_sig_rx =902;
24070: waveform_sig_rx =589;
24071: waveform_sig_rx =809;
24072: waveform_sig_rx =690;
24073: waveform_sig_rx =728;
24074: waveform_sig_rx =656;
24075: waveform_sig_rx =667;
24076: waveform_sig_rx =848;
24077: waveform_sig_rx =467;
24078: waveform_sig_rx =820;
24079: waveform_sig_rx =742;
24080: waveform_sig_rx =473;
24081: waveform_sig_rx =809;
24082: waveform_sig_rx =715;
24083: waveform_sig_rx =486;
24084: waveform_sig_rx =703;
24085: waveform_sig_rx =784;
24086: waveform_sig_rx =458;
24087: waveform_sig_rx =617;
24088: waveform_sig_rx =834;
24089: waveform_sig_rx =438;
24090: waveform_sig_rx =525;
24091: waveform_sig_rx =840;
24092: waveform_sig_rx =447;
24093: waveform_sig_rx =562;
24094: waveform_sig_rx =607;
24095: waveform_sig_rx =656;
24096: waveform_sig_rx =460;
24097: waveform_sig_rx =573;
24098: waveform_sig_rx =706;
24099: waveform_sig_rx =428;
24100: waveform_sig_rx =494;
24101: waveform_sig_rx =732;
24102: waveform_sig_rx =453;
24103: waveform_sig_rx =392;
24104: waveform_sig_rx =718;
24105: waveform_sig_rx =495;
24106: waveform_sig_rx =362;
24107: waveform_sig_rx =646;
24108: waveform_sig_rx =558;
24109: waveform_sig_rx =340;
24110: waveform_sig_rx =616;
24111: waveform_sig_rx =337;
24112: waveform_sig_rx =578;
24113: waveform_sig_rx =399;
24114: waveform_sig_rx =501;
24115: waveform_sig_rx =399;
24116: waveform_sig_rx =403;
24117: waveform_sig_rx =576;
24118: waveform_sig_rx =225;
24119: waveform_sig_rx =556;
24120: waveform_sig_rx =481;
24121: waveform_sig_rx =219;
24122: waveform_sig_rx =529;
24123: waveform_sig_rx =504;
24124: waveform_sig_rx =156;
24125: waveform_sig_rx =506;
24126: waveform_sig_rx =528;
24127: waveform_sig_rx =131;
24128: waveform_sig_rx =457;
24129: waveform_sig_rx =497;
24130: waveform_sig_rx =177;
24131: waveform_sig_rx =332;
24132: waveform_sig_rx =464;
24133: waveform_sig_rx =236;
24134: waveform_sig_rx =287;
24135: waveform_sig_rx =324;
24136: waveform_sig_rx =450;
24137: waveform_sig_rx =118;
24138: waveform_sig_rx =328;
24139: waveform_sig_rx =432;
24140: waveform_sig_rx =91;
24141: waveform_sig_rx =263;
24142: waveform_sig_rx =448;
24143: waveform_sig_rx =145;
24144: waveform_sig_rx =162;
24145: waveform_sig_rx =418;
24146: waveform_sig_rx =204;
24147: waveform_sig_rx =94;
24148: waveform_sig_rx =342;
24149: waveform_sig_rx =272;
24150: waveform_sig_rx =86;
24151: waveform_sig_rx =301;
24152: waveform_sig_rx =78;
24153: waveform_sig_rx =295;
24154: waveform_sig_rx =80;
24155: waveform_sig_rx =257;
24156: waveform_sig_rx =57;
24157: waveform_sig_rx =128;
24158: waveform_sig_rx =292;
24159: waveform_sig_rx =-124;
24160: waveform_sig_rx =258;
24161: waveform_sig_rx =196;
24162: waveform_sig_rx =-151;
24163: waveform_sig_rx =302;
24164: waveform_sig_rx =161;
24165: waveform_sig_rx =-192;
24166: waveform_sig_rx =286;
24167: waveform_sig_rx =120;
24168: waveform_sig_rx =-130;
24169: waveform_sig_rx =187;
24170: waveform_sig_rx =116;
24171: waveform_sig_rx =-35;
24172: waveform_sig_rx =-8;
24173: waveform_sig_rx =186;
24174: waveform_sig_rx =1;
24175: waveform_sig_rx =-77;
24176: waveform_sig_rx =99;
24177: waveform_sig_rx =120;
24178: waveform_sig_rx =-203;
24179: waveform_sig_rx =90;
24180: waveform_sig_rx =109;
24181: waveform_sig_rx =-181;
24182: waveform_sig_rx =-36;
24183: waveform_sig_rx =133;
24184: waveform_sig_rx =-165;
24185: waveform_sig_rx =-142;
24186: waveform_sig_rx =99;
24187: waveform_sig_rx =-134;
24188: waveform_sig_rx =-185;
24189: waveform_sig_rx =-16;
24190: waveform_sig_rx =-27;
24191: waveform_sig_rx =-228;
24192: waveform_sig_rx =-47;
24193: waveform_sig_rx =-163;
24194: waveform_sig_rx =-68;
24195: waveform_sig_rx =-200;
24196: waveform_sig_rx =3;
24197: waveform_sig_rx =-301;
24198: waveform_sig_rx =-91;
24199: waveform_sig_rx =-43;
24200: waveform_sig_rx =-440;
24201: waveform_sig_rx =39;
24202: waveform_sig_rx =-201;
24203: waveform_sig_rx =-378;
24204: waveform_sig_rx =20;
24205: waveform_sig_rx =-196;
24206: waveform_sig_rx =-417;
24207: waveform_sig_rx =-59;
24208: waveform_sig_rx =-168;
24209: waveform_sig_rx =-396;
24210: waveform_sig_rx =-152;
24211: waveform_sig_rx =-165;
24212: waveform_sig_rx =-363;
24213: waveform_sig_rx =-319;
24214: waveform_sig_rx =-118;
24215: waveform_sig_rx =-334;
24216: waveform_sig_rx =-413;
24217: waveform_sig_rx =-193;
24218: waveform_sig_rx =-216;
24219: waveform_sig_rx =-532;
24220: waveform_sig_rx =-188;
24221: waveform_sig_rx =-262;
24222: waveform_sig_rx =-504;
24223: waveform_sig_rx =-292;
24224: waveform_sig_rx =-226;
24225: waveform_sig_rx =-430;
24226: waveform_sig_rx =-444;
24227: waveform_sig_rx =-235;
24228: waveform_sig_rx =-371;
24229: waveform_sig_rx =-536;
24230: waveform_sig_rx =-276;
24231: waveform_sig_rx =-295;
24232: waveform_sig_rx =-602;
24233: waveform_sig_rx =-272;
24234: waveform_sig_rx =-490;
24235: waveform_sig_rx =-402;
24236: waveform_sig_rx =-447;
24237: waveform_sig_rx =-359;
24238: waveform_sig_rx =-619;
24239: waveform_sig_rx =-333;
24240: waveform_sig_rx =-400;
24241: waveform_sig_rx =-670;
24242: waveform_sig_rx =-252;
24243: waveform_sig_rx =-514;
24244: waveform_sig_rx =-623;
24245: waveform_sig_rx =-326;
24246: waveform_sig_rx =-490;
24247: waveform_sig_rx =-697;
24248: waveform_sig_rx =-365;
24249: waveform_sig_rx =-470;
24250: waveform_sig_rx =-684;
24251: waveform_sig_rx =-452;
24252: waveform_sig_rx =-446;
24253: waveform_sig_rx =-662;
24254: waveform_sig_rx =-627;
24255: waveform_sig_rx =-355;
24256: waveform_sig_rx =-649;
24257: waveform_sig_rx =-669;
24258: waveform_sig_rx =-428;
24259: waveform_sig_rx =-578;
24260: waveform_sig_rx =-754;
24261: waveform_sig_rx =-451;
24262: waveform_sig_rx =-595;
24263: waveform_sig_rx =-693;
24264: waveform_sig_rx =-624;
24265: waveform_sig_rx =-478;
24266: waveform_sig_rx =-679;
24267: waveform_sig_rx =-780;
24268: waveform_sig_rx =-429;
24269: waveform_sig_rx =-683;
24270: waveform_sig_rx =-831;
24271: waveform_sig_rx =-493;
24272: waveform_sig_rx =-640;
24273: waveform_sig_rx =-839;
24274: waveform_sig_rx =-538;
24275: waveform_sig_rx =-805;
24276: waveform_sig_rx =-625;
24277: waveform_sig_rx =-732;
24278: waveform_sig_rx =-671;
24279: waveform_sig_rx =-834;
24280: waveform_sig_rx =-609;
24281: waveform_sig_rx =-692;
24282: waveform_sig_rx =-888;
24283: waveform_sig_rx =-565;
24284: waveform_sig_rx =-771;
24285: waveform_sig_rx =-873;
24286: waveform_sig_rx =-628;
24287: waveform_sig_rx =-730;
24288: waveform_sig_rx =-967;
24289: waveform_sig_rx =-641;
24290: waveform_sig_rx =-696;
24291: waveform_sig_rx =-968;
24292: waveform_sig_rx =-699;
24293: waveform_sig_rx =-668;
24294: waveform_sig_rx =-994;
24295: waveform_sig_rx =-822;
24296: waveform_sig_rx =-600;
24297: waveform_sig_rx =-958;
24298: waveform_sig_rx =-854;
24299: waveform_sig_rx =-711;
24300: waveform_sig_rx =-820;
24301: waveform_sig_rx =-963;
24302: waveform_sig_rx =-768;
24303: waveform_sig_rx =-758;
24304: waveform_sig_rx =-982;
24305: waveform_sig_rx =-871;
24306: waveform_sig_rx =-639;
24307: waveform_sig_rx =-990;
24308: waveform_sig_rx =-951;
24309: waveform_sig_rx =-655;
24310: waveform_sig_rx =-980;
24311: waveform_sig_rx =-1010;
24312: waveform_sig_rx =-747;
24313: waveform_sig_rx =-895;
24314: waveform_sig_rx =-1027;
24315: waveform_sig_rx =-771;
24316: waveform_sig_rx =-1029;
24317: waveform_sig_rx =-832;
24318: waveform_sig_rx =-987;
24319: waveform_sig_rx =-870;
24320: waveform_sig_rx =-1048;
24321: waveform_sig_rx =-864;
24322: waveform_sig_rx =-920;
24323: waveform_sig_rx =-1106;
24324: waveform_sig_rx =-831;
24325: waveform_sig_rx =-942;
24326: waveform_sig_rx =-1136;
24327: waveform_sig_rx =-800;
24328: waveform_sig_rx =-901;
24329: waveform_sig_rx =-1272;
24330: waveform_sig_rx =-761;
24331: waveform_sig_rx =-962;
24332: waveform_sig_rx =-1221;
24333: waveform_sig_rx =-809;
24334: waveform_sig_rx =-946;
24335: waveform_sig_rx =-1160;
24336: waveform_sig_rx =-967;
24337: waveform_sig_rx =-878;
24338: waveform_sig_rx =-1101;
24339: waveform_sig_rx =-1057;
24340: waveform_sig_rx =-925;
24341: waveform_sig_rx =-973;
24342: waveform_sig_rx =-1180;
24343: waveform_sig_rx =-932;
24344: waveform_sig_rx =-936;
24345: waveform_sig_rx =-1185;
24346: waveform_sig_rx =-1044;
24347: waveform_sig_rx =-822;
24348: waveform_sig_rx =-1227;
24349: waveform_sig_rx =-1085;
24350: waveform_sig_rx =-821;
24351: waveform_sig_rx =-1206;
24352: waveform_sig_rx =-1090;
24353: waveform_sig_rx =-925;
24354: waveform_sig_rx =-1074;
24355: waveform_sig_rx =-1118;
24356: waveform_sig_rx =-1013;
24357: waveform_sig_rx =-1152;
24358: waveform_sig_rx =-977;
24359: waveform_sig_rx =-1181;
24360: waveform_sig_rx =-968;
24361: waveform_sig_rx =-1231;
24362: waveform_sig_rx =-1019;
24363: waveform_sig_rx =-1026;
24364: waveform_sig_rx =-1297;
24365: waveform_sig_rx =-896;
24366: waveform_sig_rx =-1089;
24367: waveform_sig_rx =-1314;
24368: waveform_sig_rx =-855;
24369: waveform_sig_rx =-1111;
24370: waveform_sig_rx =-1366;
24371: waveform_sig_rx =-837;
24372: waveform_sig_rx =-1183;
24373: waveform_sig_rx =-1300;
24374: waveform_sig_rx =-952;
24375: waveform_sig_rx =-1113;
24376: waveform_sig_rx =-1248;
24377: waveform_sig_rx =-1106;
24378: waveform_sig_rx =-1016;
24379: waveform_sig_rx =-1200;
24380: waveform_sig_rx =-1218;
24381: waveform_sig_rx =-1025;
24382: waveform_sig_rx =-1084;
24383: waveform_sig_rx =-1320;
24384: waveform_sig_rx =-992;
24385: waveform_sig_rx =-1066;
24386: waveform_sig_rx =-1345;
24387: waveform_sig_rx =-1056;
24388: waveform_sig_rx =-983;
24389: waveform_sig_rx =-1322;
24390: waveform_sig_rx =-1120;
24391: waveform_sig_rx =-1006;
24392: waveform_sig_rx =-1259;
24393: waveform_sig_rx =-1184;
24394: waveform_sig_rx =-1059;
24395: waveform_sig_rx =-1121;
24396: waveform_sig_rx =-1244;
24397: waveform_sig_rx =-1115;
24398: waveform_sig_rx =-1177;
24399: waveform_sig_rx =-1105;
24400: waveform_sig_rx =-1241;
24401: waveform_sig_rx =-1011;
24402: waveform_sig_rx =-1359;
24403: waveform_sig_rx =-989;
24404: waveform_sig_rx =-1138;
24405: waveform_sig_rx =-1367;
24406: waveform_sig_rx =-906;
24407: waveform_sig_rx =-1251;
24408: waveform_sig_rx =-1322;
24409: waveform_sig_rx =-915;
24410: waveform_sig_rx =-1244;
24411: waveform_sig_rx =-1336;
24412: waveform_sig_rx =-913;
24413: waveform_sig_rx =-1227;
24414: waveform_sig_rx =-1272;
24415: waveform_sig_rx =-1036;
24416: waveform_sig_rx =-1124;
24417: waveform_sig_rx =-1275;
24418: waveform_sig_rx =-1143;
24419: waveform_sig_rx =-1038;
24420: waveform_sig_rx =-1225;
24421: waveform_sig_rx =-1248;
24422: waveform_sig_rx =-1009;
24423: waveform_sig_rx =-1127;
24424: waveform_sig_rx =-1366;
24425: waveform_sig_rx =-939;
24426: waveform_sig_rx =-1154;
24427: waveform_sig_rx =-1301;
24428: waveform_sig_rx =-1036;
24429: waveform_sig_rx =-1096;
24430: waveform_sig_rx =-1257;
24431: waveform_sig_rx =-1172;
24432: waveform_sig_rx =-1030;
24433: waveform_sig_rx =-1182;
24434: waveform_sig_rx =-1271;
24435: waveform_sig_rx =-993;
24436: waveform_sig_rx =-1118;
24437: waveform_sig_rx =-1273;
24438: waveform_sig_rx =-1018;
24439: waveform_sig_rx =-1216;
24440: waveform_sig_rx =-1085;
24441: waveform_sig_rx =-1157;
24442: waveform_sig_rx =-1048;
24443: waveform_sig_rx =-1335;
24444: waveform_sig_rx =-929;
24445: waveform_sig_rx =-1187;
24446: waveform_sig_rx =-1302;
24447: waveform_sig_rx =-868;
24448: waveform_sig_rx =-1295;
24449: waveform_sig_rx =-1201;
24450: waveform_sig_rx =-893;
24451: waveform_sig_rx =-1236;
24452: waveform_sig_rx =-1238;
24453: waveform_sig_rx =-956;
24454: waveform_sig_rx =-1168;
24455: waveform_sig_rx =-1220;
24456: waveform_sig_rx =-1046;
24457: waveform_sig_rx =-1008;
24458: waveform_sig_rx =-1295;
24459: waveform_sig_rx =-1086;
24460: waveform_sig_rx =-950;
24461: waveform_sig_rx =-1236;
24462: waveform_sig_rx =-1168;
24463: waveform_sig_rx =-943;
24464: waveform_sig_rx =-1138;
24465: waveform_sig_rx =-1247;
24466: waveform_sig_rx =-909;
24467: waveform_sig_rx =-1118;
24468: waveform_sig_rx =-1217;
24469: waveform_sig_rx =-1004;
24470: waveform_sig_rx =-1006;
24471: waveform_sig_rx =-1169;
24472: waveform_sig_rx =-1118;
24473: waveform_sig_rx =-931;
24474: waveform_sig_rx =-1125;
24475: waveform_sig_rx =-1235;
24476: waveform_sig_rx =-848;
24477: waveform_sig_rx =-1114;
24478: waveform_sig_rx =-1175;
24479: waveform_sig_rx =-903;
24480: waveform_sig_rx =-1209;
24481: waveform_sig_rx =-955;
24482: waveform_sig_rx =-1100;
24483: waveform_sig_rx =-1000;
24484: waveform_sig_rx =-1173;
24485: waveform_sig_rx =-843;
24486: waveform_sig_rx =-1121;
24487: waveform_sig_rx =-1127;
24488: waveform_sig_rx =-844;
24489: waveform_sig_rx =-1168;
24490: waveform_sig_rx =-1088;
24491: waveform_sig_rx =-818;
24492: waveform_sig_rx =-1090;
24493: waveform_sig_rx =-1146;
24494: waveform_sig_rx =-828;
24495: waveform_sig_rx =-1051;
24496: waveform_sig_rx =-1125;
24497: waveform_sig_rx =-884;
24498: waveform_sig_rx =-881;
24499: waveform_sig_rx =-1188;
24500: waveform_sig_rx =-902;
24501: waveform_sig_rx =-837;
24502: waveform_sig_rx =-1129;
24503: waveform_sig_rx =-972;
24504: waveform_sig_rx =-837;
24505: waveform_sig_rx =-1011;
24506: waveform_sig_rx =-1061;
24507: waveform_sig_rx =-830;
24508: waveform_sig_rx =-970;
24509: waveform_sig_rx =-1057;
24510: waveform_sig_rx =-917;
24511: waveform_sig_rx =-814;
24512: waveform_sig_rx =-1088;
24513: waveform_sig_rx =-993;
24514: waveform_sig_rx =-715;
24515: waveform_sig_rx =-1081;
24516: waveform_sig_rx =-1016;
24517: waveform_sig_rx =-684;
24518: waveform_sig_rx =-1047;
24519: waveform_sig_rx =-932;
24520: waveform_sig_rx =-821;
24521: waveform_sig_rx =-1056;
24522: waveform_sig_rx =-740;
24523: waveform_sig_rx =-971;
24524: waveform_sig_rx =-809;
24525: waveform_sig_rx =-1009;
24526: waveform_sig_rx =-745;
24527: waveform_sig_rx =-896;
24528: waveform_sig_rx =-968;
24529: waveform_sig_rx =-672;
24530: waveform_sig_rx =-952;
24531: waveform_sig_rx =-949;
24532: waveform_sig_rx =-640;
24533: waveform_sig_rx =-921;
24534: waveform_sig_rx =-981;
24535: waveform_sig_rx =-627;
24536: waveform_sig_rx =-859;
24537: waveform_sig_rx =-968;
24538: waveform_sig_rx =-653;
24539: waveform_sig_rx =-735;
24540: waveform_sig_rx =-1034;
24541: waveform_sig_rx =-650;
24542: waveform_sig_rx =-722;
24543: waveform_sig_rx =-914;
24544: waveform_sig_rx =-736;
24545: waveform_sig_rx =-701;
24546: waveform_sig_rx =-771;
24547: waveform_sig_rx =-887;
24548: waveform_sig_rx =-646;
24549: waveform_sig_rx =-685;
24550: waveform_sig_rx =-933;
24551: waveform_sig_rx =-647;
24552: waveform_sig_rx =-596;
24553: waveform_sig_rx =-959;
24554: waveform_sig_rx =-684;
24555: waveform_sig_rx =-567;
24556: waveform_sig_rx =-874;
24557: waveform_sig_rx =-753;
24558: waveform_sig_rx =-548;
24559: waveform_sig_rx =-781;
24560: waveform_sig_rx =-727;
24561: waveform_sig_rx =-660;
24562: waveform_sig_rx =-761;
24563: waveform_sig_rx =-563;
24564: waveform_sig_rx =-772;
24565: waveform_sig_rx =-544;
24566: waveform_sig_rx =-822;
24567: waveform_sig_rx =-486;
24568: waveform_sig_rx =-727;
24569: waveform_sig_rx =-765;
24570: waveform_sig_rx =-424;
24571: waveform_sig_rx =-744;
24572: waveform_sig_rx =-723;
24573: waveform_sig_rx =-407;
24574: waveform_sig_rx =-697;
24575: waveform_sig_rx =-771;
24576: waveform_sig_rx =-345;
24577: waveform_sig_rx =-698;
24578: waveform_sig_rx =-735;
24579: waveform_sig_rx =-374;
24580: waveform_sig_rx =-594;
24581: waveform_sig_rx =-737;
24582: waveform_sig_rx =-428;
24583: waveform_sig_rx =-565;
24584: waveform_sig_rx =-583;
24585: waveform_sig_rx =-609;
24586: waveform_sig_rx =-433;
24587: waveform_sig_rx =-496;
24588: waveform_sig_rx =-731;
24589: waveform_sig_rx =-283;
24590: waveform_sig_rx =-530;
24591: waveform_sig_rx =-675;
24592: waveform_sig_rx =-317;
24593: waveform_sig_rx =-430;
24594: waveform_sig_rx =-622;
24595: waveform_sig_rx =-442;
24596: waveform_sig_rx =-350;
24597: waveform_sig_rx =-575;
24598: waveform_sig_rx =-517;
24599: waveform_sig_rx =-265;
24600: waveform_sig_rx =-533;
24601: waveform_sig_rx =-441;
24602: waveform_sig_rx =-405;
24603: waveform_sig_rx =-463;
24604: waveform_sig_rx =-322;
24605: waveform_sig_rx =-522;
24606: waveform_sig_rx =-268;
24607: waveform_sig_rx =-607;
24608: waveform_sig_rx =-207;
24609: waveform_sig_rx =-434;
24610: waveform_sig_rx =-532;
24611: waveform_sig_rx =-106;
24612: waveform_sig_rx =-530;
24613: waveform_sig_rx =-452;
24614: waveform_sig_rx =-64;
24615: waveform_sig_rx =-531;
24616: waveform_sig_rx =-417;
24617: waveform_sig_rx =-102;
24618: waveform_sig_rx =-461;
24619: waveform_sig_rx =-350;
24620: waveform_sig_rx =-177;
24621: waveform_sig_rx =-293;
24622: waveform_sig_rx =-424;
24623: waveform_sig_rx =-209;
24624: waveform_sig_rx =-195;
24625: waveform_sig_rx =-344;
24626: waveform_sig_rx =-349;
24627: waveform_sig_rx =-55;
24628: waveform_sig_rx =-308;
24629: waveform_sig_rx =-394;
24630: waveform_sig_rx =-12;
24631: waveform_sig_rx =-302;
24632: waveform_sig_rx =-353;
24633: waveform_sig_rx =-80;
24634: waveform_sig_rx =-159;
24635: waveform_sig_rx =-332;
24636: waveform_sig_rx =-168;
24637: waveform_sig_rx =-57;
24638: waveform_sig_rx =-302;
24639: waveform_sig_rx =-229;
24640: waveform_sig_rx =-7;
24641: waveform_sig_rx =-232;
24642: waveform_sig_rx =-202;
24643: waveform_sig_rx =-92;
24644: waveform_sig_rx =-162;
24645: waveform_sig_rx =-90;
24646: waveform_sig_rx =-146;
24647: waveform_sig_rx =-11;
24648: waveform_sig_rx =-324;
24649: waveform_sig_rx =168;
24650: waveform_sig_rx =-231;
24651: waveform_sig_rx =-182;
24652: waveform_sig_rx =186;
24653: waveform_sig_rx =-301;
24654: waveform_sig_rx =-45;
24655: waveform_sig_rx =147;
24656: waveform_sig_rx =-236;
24657: waveform_sig_rx =-65;
24658: waveform_sig_rx =131;
24659: waveform_sig_rx =-118;
24660: waveform_sig_rx =-71;
24661: waveform_sig_rx =94;
24662: waveform_sig_rx =61;
24663: waveform_sig_rx =-189;
24664: waveform_sig_rx =114;
24665: waveform_sig_rx =107;
24666: waveform_sig_rx =-113;
24667: waveform_sig_rx =3;
24668: waveform_sig_rx =196;
24669: waveform_sig_rx =-44;
24670: waveform_sig_rx =-56;
24671: waveform_sig_rx =254;
24672: waveform_sig_rx =-4;
24673: waveform_sig_rx =-41;
24674: waveform_sig_rx =208;
24675: waveform_sig_rx =113;
24676: waveform_sig_rx =-39;
24677: waveform_sig_rx =134;
24678: waveform_sig_rx =221;
24679: waveform_sig_rx =41;
24680: waveform_sig_rx =22;
24681: waveform_sig_rx =351;
24682: waveform_sig_rx =40;
24683: waveform_sig_rx =61;
24684: waveform_sig_rx =254;
24685: waveform_sig_rx =56;
24686: waveform_sig_rx =208;
24687: waveform_sig_rx =181;
24688: waveform_sig_rx =182;
24689: waveform_sig_rx =57;
24690: waveform_sig_rx =428;
24691: waveform_sig_rx =1;
24692: waveform_sig_rx =200;
24693: waveform_sig_rx =378;
24694: waveform_sig_rx =49;
24695: waveform_sig_rx =229;
24696: waveform_sig_rx =408;
24697: waveform_sig_rx =128;
24698: waveform_sig_rx =185;
24699: waveform_sig_rx =476;
24700: waveform_sig_rx =167;
24701: waveform_sig_rx =220;
24702: waveform_sig_rx =387;
24703: waveform_sig_rx =319;
24704: waveform_sig_rx =102;
24705: waveform_sig_rx =411;
24706: waveform_sig_rx =389;
24707: waveform_sig_rx =158;
24708: waveform_sig_rx =309;
24709: waveform_sig_rx =491;
24710: waveform_sig_rx =212;
24711: waveform_sig_rx =298;
24712: waveform_sig_rx =492;
24713: waveform_sig_rx =300;
24714: waveform_sig_rx =282;
24715: waveform_sig_rx =427;
24716: waveform_sig_rx =483;
24717: waveform_sig_rx =197;
24718: waveform_sig_rx =408;
24719: waveform_sig_rx =564;
24720: waveform_sig_rx =225;
24721: waveform_sig_rx =365;
24722: waveform_sig_rx =621;
24723: waveform_sig_rx =265;
24724: waveform_sig_rx =440;
24725: waveform_sig_rx =470;
24726: waveform_sig_rx =360;
24727: waveform_sig_rx =548;
24728: waveform_sig_rx =415;
24729: waveform_sig_rx =481;
24730: waveform_sig_rx =361;
24731: waveform_sig_rx =645;
24732: waveform_sig_rx =338;
24733: waveform_sig_rx =484;
24734: waveform_sig_rx =628;
24735: waveform_sig_rx =365;
24736: waveform_sig_rx =476;
24737: waveform_sig_rx =696;
24738: waveform_sig_rx =408;
24739: waveform_sig_rx =419;
24740: waveform_sig_rx =776;
24741: waveform_sig_rx =396;
24742: waveform_sig_rx =457;
24743: waveform_sig_rx =719;
24744: waveform_sig_rx =551;
24745: waveform_sig_rx =366;
24746: waveform_sig_rx =735;
24747: waveform_sig_rx =607;
24748: waveform_sig_rx =436;
24749: waveform_sig_rx =614;
24750: waveform_sig_rx =720;
24751: waveform_sig_rx =490;
24752: waveform_sig_rx =567;
24753: waveform_sig_rx =731;
24754: waveform_sig_rx =601;
24755: waveform_sig_rx =502;
24756: waveform_sig_rx =719;
24757: waveform_sig_rx =761;
24758: waveform_sig_rx =407;
24759: waveform_sig_rx =758;
24760: waveform_sig_rx =803;
24761: waveform_sig_rx =459;
24762: waveform_sig_rx =707;
24763: waveform_sig_rx =834;
24764: waveform_sig_rx =548;
24765: waveform_sig_rx =715;
24766: waveform_sig_rx =677;
24767: waveform_sig_rx =680;
24768: waveform_sig_rx =757;
24769: waveform_sig_rx =637;
24770: waveform_sig_rx =774;
24771: waveform_sig_rx =593;
24772: waveform_sig_rx =899;
24773: waveform_sig_rx =601;
24774: waveform_sig_rx =704;
24775: waveform_sig_rx =902;
24776: waveform_sig_rx =608;
24777: waveform_sig_rx =709;
24778: waveform_sig_rx =981;
24779: waveform_sig_rx =617;
24780: waveform_sig_rx =677;
24781: waveform_sig_rx =1056;
24782: waveform_sig_rx =587;
24783: waveform_sig_rx =721;
24784: waveform_sig_rx =971;
24785: waveform_sig_rx =731;
24786: waveform_sig_rx =646;
24787: waveform_sig_rx =961;
24788: waveform_sig_rx =815;
24789: waveform_sig_rx =740;
24790: waveform_sig_rx =821;
24791: waveform_sig_rx =959;
24792: waveform_sig_rx =741;
24793: waveform_sig_rx =772;
24794: waveform_sig_rx =1003;
24795: waveform_sig_rx =825;
24796: waveform_sig_rx =715;
24797: waveform_sig_rx =1006;
24798: waveform_sig_rx =927;
24799: waveform_sig_rx =651;
24800: waveform_sig_rx =1022;
24801: waveform_sig_rx =951;
24802: waveform_sig_rx =724;
24803: waveform_sig_rx =929;
24804: waveform_sig_rx =1016;
24805: waveform_sig_rx =809;
24806: waveform_sig_rx =920;
24807: waveform_sig_rx =873;
24808: waveform_sig_rx =943;
24809: waveform_sig_rx =917;
24810: waveform_sig_rx =908;
24811: waveform_sig_rx =985;
24812: waveform_sig_rx =763;
24813: waveform_sig_rx =1155;
24814: waveform_sig_rx =793;
24815: waveform_sig_rx =904;
24816: waveform_sig_rx =1164;
24817: waveform_sig_rx =752;
24818: waveform_sig_rx =938;
24819: waveform_sig_rx =1194;
24820: waveform_sig_rx =746;
24821: waveform_sig_rx =924;
24822: waveform_sig_rx =1202;
24823: waveform_sig_rx =759;
24824: waveform_sig_rx =977;
24825: waveform_sig_rx =1103;
24826: waveform_sig_rx =916;
24827: waveform_sig_rx =861;
24828: waveform_sig_rx =1111;
24829: waveform_sig_rx =1014;
24830: waveform_sig_rx =912;
24831: waveform_sig_rx =959;
24832: waveform_sig_rx =1173;
24833: waveform_sig_rx =875;
24834: waveform_sig_rx =943;
24835: waveform_sig_rx =1207;
24836: waveform_sig_rx =912;
24837: waveform_sig_rx =898;
24838: waveform_sig_rx =1211;
24839: waveform_sig_rx =1007;
24840: waveform_sig_rx =882;
24841: waveform_sig_rx =1167;
24842: waveform_sig_rx =1080;
24843: waveform_sig_rx =937;
24844: waveform_sig_rx =1029;
24845: waveform_sig_rx =1190;
24846: waveform_sig_rx =961;
24847: waveform_sig_rx =1035;
24848: waveform_sig_rx =1096;
24849: waveform_sig_rx =1054;
24850: waveform_sig_rx =1049;
24851: waveform_sig_rx =1119;
24852: waveform_sig_rx =1072;
24853: waveform_sig_rx =962;
24854: waveform_sig_rx =1324;
24855: waveform_sig_rx =852;
24856: waveform_sig_rx =1117;
24857: waveform_sig_rx =1250;
24858: waveform_sig_rx =861;
24859: waveform_sig_rx =1135;
24860: waveform_sig_rx =1282;
24861: waveform_sig_rx =851;
24862: waveform_sig_rx =1128;
24863: waveform_sig_rx =1288;
24864: waveform_sig_rx =871;
24865: waveform_sig_rx =1153;
24866: waveform_sig_rx =1165;
24867: waveform_sig_rx =1065;
24868: waveform_sig_rx =987;
24869: waveform_sig_rx =1206;
24870: waveform_sig_rx =1160;
24871: waveform_sig_rx =959;
24872: waveform_sig_rx =1126;
24873: waveform_sig_rx =1303;
24874: waveform_sig_rx =918;
24875: waveform_sig_rx =1150;
24876: waveform_sig_rx =1302;
24877: waveform_sig_rx =1004;
24878: waveform_sig_rx =1072;
24879: waveform_sig_rx =1237;
24880: waveform_sig_rx =1120;
24881: waveform_sig_rx =977;
24882: waveform_sig_rx =1222;
24883: waveform_sig_rx =1226;
24884: waveform_sig_rx =989;
24885: waveform_sig_rx =1116;
24886: waveform_sig_rx =1325;
24887: waveform_sig_rx =963;
24888: waveform_sig_rx =1140;
24889: waveform_sig_rx =1161;
24890: waveform_sig_rx =1090;
24891: waveform_sig_rx =1154;
24892: waveform_sig_rx =1169;
24893: waveform_sig_rx =1096;
24894: waveform_sig_rx =1063;
24895: waveform_sig_rx =1337;
24896: waveform_sig_rx =909;
24897: waveform_sig_rx =1225;
24898: waveform_sig_rx =1267;
24899: waveform_sig_rx =929;
24900: waveform_sig_rx =1249;
24901: waveform_sig_rx =1265;
24902: waveform_sig_rx =935;
24903: waveform_sig_rx =1189;
24904: waveform_sig_rx =1264;
24905: waveform_sig_rx =985;
24906: waveform_sig_rx =1150;
24907: waveform_sig_rx =1243;
24908: waveform_sig_rx =1151;
24909: waveform_sig_rx =942;
24910: waveform_sig_rx =1331;
24911: waveform_sig_rx =1186;
24912: waveform_sig_rx =972;
24913: waveform_sig_rx =1237;
24914: waveform_sig_rx =1264;
24915: waveform_sig_rx =980;
24916: waveform_sig_rx =1200;
24917: waveform_sig_rx =1246;
24918: waveform_sig_rx =1085;
24919: waveform_sig_rx =1083;
24920: waveform_sig_rx =1262;
24921: waveform_sig_rx =1191;
24922: waveform_sig_rx =972;
24923: waveform_sig_rx =1246;
24924: waveform_sig_rx =1237;
24925: waveform_sig_rx =954;
24926: waveform_sig_rx =1174;
24927: waveform_sig_rx =1335;
24928: waveform_sig_rx =941;
24929: waveform_sig_rx =1229;
24930: waveform_sig_rx =1118;
24931: waveform_sig_rx =1094;
24932: waveform_sig_rx =1179;
24933: waveform_sig_rx =1143;
24934: waveform_sig_rx =1093;
24935: waveform_sig_rx =1122;
24936: waveform_sig_rx =1300;
24937: waveform_sig_rx =906;
24938: waveform_sig_rx =1252;
24939: waveform_sig_rx =1198;
24940: waveform_sig_rx =968;
24941: waveform_sig_rx =1215;
24942: waveform_sig_rx =1247;
24943: waveform_sig_rx =988;
24944: waveform_sig_rx =1112;
24945: waveform_sig_rx =1325;
24946: waveform_sig_rx =957;
24947: waveform_sig_rx =1106;
24948: waveform_sig_rx =1308;
24949: waveform_sig_rx =1051;
24950: waveform_sig_rx =978;
24951: waveform_sig_rx =1341;
24952: waveform_sig_rx =1048;
24953: waveform_sig_rx =1021;
24954: waveform_sig_rx =1160;
24955: waveform_sig_rx =1199;
24956: waveform_sig_rx =968;
24957: waveform_sig_rx =1117;
24958: waveform_sig_rx =1233;
24959: waveform_sig_rx =1018;
24960: waveform_sig_rx =1020;
24961: waveform_sig_rx =1222;
24962: waveform_sig_rx =1132;
24963: waveform_sig_rx =894;
24964: waveform_sig_rx =1235;
24965: waveform_sig_rx =1174;
24966: waveform_sig_rx =861;
24967: waveform_sig_rx =1195;
24968: waveform_sig_rx =1221;
24969: waveform_sig_rx =872;
24970: waveform_sig_rx =1245;
24971: waveform_sig_rx =954;
24972: waveform_sig_rx =1113;
24973: waveform_sig_rx =1107;
24974: waveform_sig_rx =1040;
24975: waveform_sig_rx =1086;
24976: waveform_sig_rx =975;
24977: waveform_sig_rx =1230;
24978: waveform_sig_rx =863;
24979: waveform_sig_rx =1108;
24980: waveform_sig_rx =1167;
24981: waveform_sig_rx =864;
24982: waveform_sig_rx =1111;
24983: waveform_sig_rx =1208;
24984: waveform_sig_rx =827;
24985: waveform_sig_rx =1075;
24986: waveform_sig_rx =1230;
24987: waveform_sig_rx =839;
24988: waveform_sig_rx =1033;
24989: waveform_sig_rx =1198;
24990: waveform_sig_rx =895;
24991: waveform_sig_rx =892;
24992: waveform_sig_rx =1223;
24993: waveform_sig_rx =906;
24994: waveform_sig_rx =950;
24995: waveform_sig_rx =1013;
24996: waveform_sig_rx =1081;
24997: waveform_sig_rx =875;
24998: waveform_sig_rx =948;
24999: waveform_sig_rx =1148;
25000: waveform_sig_rx =890;
25001: waveform_sig_rx =876;
25002: waveform_sig_rx =1182;
25003: waveform_sig_rx =933;
25004: waveform_sig_rx =798;
25005: waveform_sig_rx =1158;
25006: waveform_sig_rx =971;
25007: waveform_sig_rx =790;
25008: waveform_sig_rx =1059;
25009: waveform_sig_rx =1026;
25010: waveform_sig_rx =810;
25011: waveform_sig_rx =1044;
25012: waveform_sig_rx =808;
25013: waveform_sig_rx =1030;
25014: waveform_sig_rx =885;
25015: waveform_sig_rx =953;
25016: waveform_sig_rx =941;
25017: waveform_sig_rx =814;
25018: waveform_sig_rx =1125;
25019: waveform_sig_rx =695;
25020: waveform_sig_rx =961;
25021: waveform_sig_rx =1046;
25022: waveform_sig_rx =639;
25023: waveform_sig_rx =1004;
25024: waveform_sig_rx =1048;
25025: waveform_sig_rx =630;
25026: waveform_sig_rx =958;
25027: waveform_sig_rx =1044;
25028: waveform_sig_rx =636;
25029: waveform_sig_rx =913;
25030: waveform_sig_rx =998;
25031: waveform_sig_rx =710;
25032: waveform_sig_rx =805;
25033: waveform_sig_rx =996;
25034: waveform_sig_rx =754;
25035: waveform_sig_rx =826;
25036: waveform_sig_rx =813;
25037: waveform_sig_rx =993;
25038: waveform_sig_rx =668;
25039: waveform_sig_rx =793;
25040: waveform_sig_rx =1019;
25041: waveform_sig_rx =603;
25042: waveform_sig_rx =771;
25043: waveform_sig_rx =986;
25044: waveform_sig_rx =691;
25045: waveform_sig_rx =705;
25046: waveform_sig_rx =909;
25047: waveform_sig_rx =763;
25048: waveform_sig_rx =634;
25049: waveform_sig_rx =827;
25050: waveform_sig_rx =864;
25051: waveform_sig_rx =592;
25052: waveform_sig_rx =837;
25053: waveform_sig_rx =626;
25054: waveform_sig_rx =809;
25055: waveform_sig_rx =683;
25056: waveform_sig_rx =786;
25057: waveform_sig_rx =675;
25058: waveform_sig_rx =633;
25059: waveform_sig_rx =931;
25060: waveform_sig_rx =437;
25061: waveform_sig_rx =807;
25062: waveform_sig_rx =832;
25063: waveform_sig_rx =387;
25064: waveform_sig_rx =859;
25065: waveform_sig_rx =781;
25066: waveform_sig_rx =368;
25067: waveform_sig_rx =822;
25068: waveform_sig_rx =720;
25069: waveform_sig_rx =449;
25070: waveform_sig_rx =738;
25071: waveform_sig_rx =691;
25072: waveform_sig_rx =565;
25073: waveform_sig_rx =534;
25074: waveform_sig_rx =760;
25075: waveform_sig_rx =590;
25076: waveform_sig_rx =480;
25077: waveform_sig_rx =631;
25078: waveform_sig_rx =727;
25079: waveform_sig_rx =364;
25080: waveform_sig_rx =650;
25081: waveform_sig_rx =711;
25082: waveform_sig_rx =388;
25083: waveform_sig_rx =568;
25084: waveform_sig_rx =684;
25085: waveform_sig_rx =470;
25086: waveform_sig_rx =434;
25087: waveform_sig_rx =630;
25088: waveform_sig_rx =525;
25089: waveform_sig_rx =361;
25090: waveform_sig_rx =560;
25091: waveform_sig_rx =625;
25092: waveform_sig_rx =338;
25093: waveform_sig_rx =564;
25094: waveform_sig_rx =415;
25095: waveform_sig_rx =522;
25096: waveform_sig_rx =418;
25097: waveform_sig_rx =558;
25098: waveform_sig_rx =342;
25099: waveform_sig_rx =437;
25100: waveform_sig_rx =635;
25101: waveform_sig_rx =126;
25102: waveform_sig_rx =627;
25103: waveform_sig_rx =477;
25104: waveform_sig_rx =158;
25105: waveform_sig_rx =629;
25106: waveform_sig_rx =397;
25107: waveform_sig_rx =209;
25108: waveform_sig_rx =516;
25109: waveform_sig_rx =419;
25110: waveform_sig_rx =260;
25111: waveform_sig_rx =371;
25112: waveform_sig_rx =481;
25113: waveform_sig_rx =262;
25114: waveform_sig_rx =199;
25115: waveform_sig_rx =555;
25116: waveform_sig_rx =256;
25117: waveform_sig_rx =223;
25118: waveform_sig_rx =394;
25119: waveform_sig_rx =422;
25120: waveform_sig_rx =104;
25121: waveform_sig_rx =382;
25122: waveform_sig_rx =407;
25123: waveform_sig_rx =114;
25124: waveform_sig_rx =295;
25125: waveform_sig_rx =370;
25126: waveform_sig_rx =204;
25127: waveform_sig_rx =150;
25128: waveform_sig_rx =342;
25129: waveform_sig_rx =278;
25130: waveform_sig_rx =50;
25131: waveform_sig_rx =293;
25132: waveform_sig_rx =342;
25133: waveform_sig_rx =-23;
25134: waveform_sig_rx =336;
25135: waveform_sig_rx =104;
25136: waveform_sig_rx =199;
25137: waveform_sig_rx =165;
25138: waveform_sig_rx =229;
25139: waveform_sig_rx =35;
25140: waveform_sig_rx =204;
25141: waveform_sig_rx =240;
25142: waveform_sig_rx =-103;
25143: waveform_sig_rx =303;
25144: waveform_sig_rx =105;
25145: waveform_sig_rx =-59;
25146: waveform_sig_rx =249;
25147: waveform_sig_rx =143;
25148: waveform_sig_rx =-84;
25149: waveform_sig_rx =176;
25150: waveform_sig_rx =179;
25151: waveform_sig_rx =-96;
25152: waveform_sig_rx =81;
25153: waveform_sig_rx =199;
25154: waveform_sig_rx =-71;
25155: waveform_sig_rx =-44;
25156: waveform_sig_rx =237;
25157: waveform_sig_rx =-72;
25158: waveform_sig_rx =-61;
25159: waveform_sig_rx =104;
25160: waveform_sig_rx =79;
25161: waveform_sig_rx =-205;
25162: waveform_sig_rx =105;
25163: waveform_sig_rx =49;
25164: waveform_sig_rx =-142;
25165: waveform_sig_rx =-48;
25166: waveform_sig_rx =70;
25167: waveform_sig_rx =-47;
25168: waveform_sig_rx =-227;
25169: waveform_sig_rx =120;
25170: waveform_sig_rx =-29;
25171: waveform_sig_rx =-306;
25172: waveform_sig_rx =102;
25173: waveform_sig_rx =-31;
25174: waveform_sig_rx =-269;
25175: waveform_sig_rx =71;
25176: waveform_sig_rx =-267;
25177: waveform_sig_rx =-22;
25178: waveform_sig_rx =-154;
25179: waveform_sig_rx =-115;
25180: waveform_sig_rx =-212;
25181: waveform_sig_rx =-142;
25182: waveform_sig_rx =-63;
25183: waveform_sig_rx =-382;
25184: waveform_sig_rx =-50;
25185: waveform_sig_rx =-137;
25186: waveform_sig_rx =-374;
25187: waveform_sig_rx =-71;
25188: waveform_sig_rx =-138;
25189: waveform_sig_rx =-426;
25190: waveform_sig_rx =-124;
25191: waveform_sig_rx =-124;
25192: waveform_sig_rx =-447;
25193: waveform_sig_rx =-176;
25194: waveform_sig_rx =-112;
25195: waveform_sig_rx =-419;
25196: waveform_sig_rx =-324;
25197: waveform_sig_rx =-69;
25198: waveform_sig_rx =-402;
25199: waveform_sig_rx =-353;
25200: waveform_sig_rx =-219;
25201: waveform_sig_rx =-256;
25202: waveform_sig_rx =-454;
25203: waveform_sig_rx =-257;
25204: waveform_sig_rx =-223;
25205: waveform_sig_rx =-441;
25206: waveform_sig_rx =-417;
25207: waveform_sig_rx =-151;
25208: waveform_sig_rx =-442;
25209: waveform_sig_rx =-512;
25210: waveform_sig_rx =-135;
25211: waveform_sig_rx =-451;
25212: waveform_sig_rx =-531;
25213: waveform_sig_rx =-215;
25214: waveform_sig_rx =-372;
25215: waveform_sig_rx =-516;
25216: waveform_sig_rx =-305;
25217: waveform_sig_rx =-541;
25218: waveform_sig_rx =-293;
25219: waveform_sig_rx =-521;
25220: waveform_sig_rx =-359;
25221: waveform_sig_rx =-527;
25222: waveform_sig_rx =-454;
25223: waveform_sig_rx =-335;
25224: waveform_sig_rx =-672;
25225: waveform_sig_rx =-351;
25226: waveform_sig_rx =-423;
25227: waveform_sig_rx =-694;
25228: waveform_sig_rx =-352;
25229: waveform_sig_rx =-415;
25230: waveform_sig_rx =-772;
25231: waveform_sig_rx =-355;
25232: waveform_sig_rx =-437;
25233: waveform_sig_rx =-773;
25234: waveform_sig_rx =-405;
25235: waveform_sig_rx =-452;
25236: waveform_sig_rx =-716;
25237: waveform_sig_rx =-569;
25238: waveform_sig_rx =-405;
25239: waveform_sig_rx =-659;
25240: waveform_sig_rx =-623;
25241: waveform_sig_rx =-515;
25242: waveform_sig_rx =-503;
25243: waveform_sig_rx =-761;
25244: waveform_sig_rx =-537;
25245: waveform_sig_rx =-464;
25246: waveform_sig_rx =-752;
25247: waveform_sig_rx =-634;
25248: waveform_sig_rx =-405;
25249: waveform_sig_rx =-783;
25250: waveform_sig_rx =-723;
25251: waveform_sig_rx =-435;
25252: waveform_sig_rx =-744;
25253: waveform_sig_rx =-722;
25254: waveform_sig_rx =-579;
25255: waveform_sig_rx =-634;
25256: waveform_sig_rx =-782;
25257: waveform_sig_rx =-628;
25258: waveform_sig_rx =-771;
25259: waveform_sig_rx =-622;
25260: waveform_sig_rx =-801;
25261: waveform_sig_rx =-594;
25262: waveform_sig_rx =-850;
25263: waveform_sig_rx =-686;
25264: waveform_sig_rx =-599;
25265: waveform_sig_rx =-995;
25266: waveform_sig_rx =-568;
25267: waveform_sig_rx =-707;
25268: waveform_sig_rx =-1000;
25269: waveform_sig_rx =-559;
25270: waveform_sig_rx =-715;
25271: waveform_sig_rx =-1033;
25272: waveform_sig_rx =-556;
25273: waveform_sig_rx =-749;
25274: waveform_sig_rx =-976;
25275: waveform_sig_rx =-643;
25276: waveform_sig_rx =-764;
25277: waveform_sig_rx =-903;
25278: waveform_sig_rx =-838;
25279: waveform_sig_rx =-680;
25280: waveform_sig_rx =-860;
25281: waveform_sig_rx =-935;
25282: waveform_sig_rx =-729;
25283: waveform_sig_rx =-745;
25284: waveform_sig_rx =-1051;
25285: waveform_sig_rx =-718;
25286: waveform_sig_rx =-752;
25287: waveform_sig_rx =-1065;
25288: waveform_sig_rx =-823;
25289: waveform_sig_rx =-706;
25290: waveform_sig_rx =-1005;
25291: waveform_sig_rx =-910;
25292: waveform_sig_rx =-756;
25293: waveform_sig_rx =-945;
25294: waveform_sig_rx =-982;
25295: waveform_sig_rx =-819;
25296: waveform_sig_rx =-802;
25297: waveform_sig_rx =-1063;
25298: waveform_sig_rx =-838;
25299: waveform_sig_rx =-942;
25300: waveform_sig_rx =-889;
25301: waveform_sig_rx =-969;
25302: waveform_sig_rx =-807;
25303: waveform_sig_rx =-1110;
25304: waveform_sig_rx =-811;
25305: waveform_sig_rx =-870;
25306: waveform_sig_rx =-1185;
25307: waveform_sig_rx =-757;
25308: waveform_sig_rx =-984;
25309: waveform_sig_rx =-1135;
25310: waveform_sig_rx =-739;
25311: waveform_sig_rx =-956;
25312: waveform_sig_rx =-1204;
25313: waveform_sig_rx =-759;
25314: waveform_sig_rx =-1001;
25315: waveform_sig_rx =-1155;
25316: waveform_sig_rx =-867;
25317: waveform_sig_rx =-971;
25318: waveform_sig_rx =-1079;
25319: waveform_sig_rx =-1062;
25320: waveform_sig_rx =-844;
25321: waveform_sig_rx =-1059;
25322: waveform_sig_rx =-1161;
25323: waveform_sig_rx =-844;
25324: waveform_sig_rx =-988;
25325: waveform_sig_rx =-1237;
25326: waveform_sig_rx =-827;
25327: waveform_sig_rx =-1024;
25328: waveform_sig_rx =-1172;
25329: waveform_sig_rx =-1013;
25330: waveform_sig_rx =-934;
25331: waveform_sig_rx =-1128;
25332: waveform_sig_rx =-1146;
25333: waveform_sig_rx =-873;
25334: waveform_sig_rx =-1088;
25335: waveform_sig_rx =-1195;
25336: waveform_sig_rx =-913;
25337: waveform_sig_rx =-1012;
25338: waveform_sig_rx =-1210;
25339: waveform_sig_rx =-966;
25340: waveform_sig_rx =-1154;
25341: waveform_sig_rx =-1029;
25342: waveform_sig_rx =-1119;
25343: waveform_sig_rx =-994;
25344: waveform_sig_rx =-1250;
25345: waveform_sig_rx =-948;
25346: waveform_sig_rx =-1049;
25347: waveform_sig_rx =-1296;
25348: waveform_sig_rx =-866;
25349: waveform_sig_rx =-1169;
25350: waveform_sig_rx =-1244;
25351: waveform_sig_rx =-905;
25352: waveform_sig_rx =-1154;
25353: waveform_sig_rx =-1274;
25354: waveform_sig_rx =-956;
25355: waveform_sig_rx =-1120;
25356: waveform_sig_rx =-1242;
25357: waveform_sig_rx =-1073;
25358: waveform_sig_rx =-1020;
25359: waveform_sig_rx =-1258;
25360: waveform_sig_rx =-1186;
25361: waveform_sig_rx =-902;
25362: waveform_sig_rx =-1261;
25363: waveform_sig_rx =-1207;
25364: waveform_sig_rx =-973;
25365: waveform_sig_rx =-1166;
25366: waveform_sig_rx =-1247;
25367: waveform_sig_rx =-1022;
25368: waveform_sig_rx =-1106;
25369: waveform_sig_rx =-1235;
25370: waveform_sig_rx =-1167;
25371: waveform_sig_rx =-972;
25372: waveform_sig_rx =-1251;
25373: waveform_sig_rx =-1242;
25374: waveform_sig_rx =-952;
25375: waveform_sig_rx =-1239;
25376: waveform_sig_rx =-1267;
25377: waveform_sig_rx =-996;
25378: waveform_sig_rx =-1132;
25379: waveform_sig_rx =-1297;
25380: waveform_sig_rx =-1031;
25381: waveform_sig_rx =-1268;
25382: waveform_sig_rx =-1088;
25383: waveform_sig_rx =-1199;
25384: waveform_sig_rx =-1103;
25385: waveform_sig_rx =-1308;
25386: waveform_sig_rx =-1023;
25387: waveform_sig_rx =-1187;
25388: waveform_sig_rx =-1316;
25389: waveform_sig_rx =-988;
25390: waveform_sig_rx =-1254;
25391: waveform_sig_rx =-1260;
25392: waveform_sig_rx =-1032;
25393: waveform_sig_rx =-1143;
25394: waveform_sig_rx =-1356;
25395: waveform_sig_rx =-1009;
25396: waveform_sig_rx =-1107;
25397: waveform_sig_rx =-1370;
25398: waveform_sig_rx =-1042;
25399: waveform_sig_rx =-1064;
25400: waveform_sig_rx =-1339;
25401: waveform_sig_rx =-1100;
25402: waveform_sig_rx =-1032;
25403: waveform_sig_rx =-1293;
25404: waveform_sig_rx =-1167;
25405: waveform_sig_rx =-1072;
25406: waveform_sig_rx =-1143;
25407: waveform_sig_rx =-1300;
25408: waveform_sig_rx =-1053;
25409: waveform_sig_rx =-1072;
25410: waveform_sig_rx =-1311;
25411: waveform_sig_rx =-1134;
25412: waveform_sig_rx =-977;
25413: waveform_sig_rx =-1305;
25414: waveform_sig_rx =-1212;
25415: waveform_sig_rx =-951;
25416: waveform_sig_rx =-1266;
25417: waveform_sig_rx =-1263;
25418: waveform_sig_rx =-974;
25419: waveform_sig_rx =-1202;
25420: waveform_sig_rx =-1238;
25421: waveform_sig_rx =-1031;
25422: waveform_sig_rx =-1310;
25423: waveform_sig_rx =-996;
25424: waveform_sig_rx =-1231;
25425: waveform_sig_rx =-1068;
25426: waveform_sig_rx =-1238;
25427: waveform_sig_rx =-1057;
25428: waveform_sig_rx =-1127;
25429: waveform_sig_rx =-1303;
25430: waveform_sig_rx =-993;
25431: waveform_sig_rx =-1153;
25432: waveform_sig_rx =-1336;
25433: waveform_sig_rx =-905;
25434: waveform_sig_rx =-1128;
25435: waveform_sig_rx =-1368;
25436: waveform_sig_rx =-839;
25437: waveform_sig_rx =-1170;
25438: waveform_sig_rx =-1280;
25439: waveform_sig_rx =-957;
25440: waveform_sig_rx =-1090;
25441: waveform_sig_rx =-1254;
25442: waveform_sig_rx =-1065;
25443: waveform_sig_rx =-998;
25444: waveform_sig_rx =-1211;
25445: waveform_sig_rx =-1145;
25446: waveform_sig_rx =-998;
25447: waveform_sig_rx =-1083;
25448: waveform_sig_rx =-1256;
25449: waveform_sig_rx =-970;
25450: waveform_sig_rx =-1043;
25451: waveform_sig_rx =-1264;
25452: waveform_sig_rx =-1056;
25453: waveform_sig_rx =-924;
25454: waveform_sig_rx =-1284;
25455: waveform_sig_rx =-1108;
25456: waveform_sig_rx =-901;
25457: waveform_sig_rx =-1228;
25458: waveform_sig_rx =-1122;
25459: waveform_sig_rx =-947;
25460: waveform_sig_rx =-1121;
25461: waveform_sig_rx =-1118;
25462: waveform_sig_rx =-1040;
25463: waveform_sig_rx =-1144;
25464: waveform_sig_rx =-946;
25465: waveform_sig_rx =-1180;
25466: waveform_sig_rx =-906;
25467: waveform_sig_rx =-1226;
25468: waveform_sig_rx =-897;
25469: waveform_sig_rx =-1002;
25470: waveform_sig_rx =-1251;
25471: waveform_sig_rx =-784;
25472: waveform_sig_rx =-1098;
25473: waveform_sig_rx =-1201;
25474: waveform_sig_rx =-733;
25475: waveform_sig_rx =-1119;
25476: waveform_sig_rx =-1197;
25477: waveform_sig_rx =-765;
25478: waveform_sig_rx =-1083;
25479: waveform_sig_rx =-1119;
25480: waveform_sig_rx =-866;
25481: waveform_sig_rx =-959;
25482: waveform_sig_rx =-1157;
25483: waveform_sig_rx =-931;
25484: waveform_sig_rx =-881;
25485: waveform_sig_rx =-1067;
25486: waveform_sig_rx =-1025;
25487: waveform_sig_rx =-855;
25488: waveform_sig_rx =-933;
25489: waveform_sig_rx =-1151;
25490: waveform_sig_rx =-780;
25491: waveform_sig_rx =-912;
25492: waveform_sig_rx =-1153;
25493: waveform_sig_rx =-807;
25494: waveform_sig_rx =-851;
25495: waveform_sig_rx =-1090;
25496: waveform_sig_rx =-904;
25497: waveform_sig_rx =-833;
25498: waveform_sig_rx =-980;
25499: waveform_sig_rx =-1004;
25500: waveform_sig_rx =-770;
25501: waveform_sig_rx =-917;
25502: waveform_sig_rx =-1018;
25503: waveform_sig_rx =-833;
25504: waveform_sig_rx =-959;
25505: waveform_sig_rx =-836;
25506: waveform_sig_rx =-953;
25507: waveform_sig_rx =-763;
25508: waveform_sig_rx =-1100;
25509: waveform_sig_rx =-665;
25510: waveform_sig_rx =-914;
25511: waveform_sig_rx =-1052;
25512: waveform_sig_rx =-589;
25513: waveform_sig_rx =-1011;
25514: waveform_sig_rx =-946;
25515: waveform_sig_rx =-573;
25516: waveform_sig_rx =-962;
25517: waveform_sig_rx =-947;
25518: waveform_sig_rx =-618;
25519: waveform_sig_rx =-937;
25520: waveform_sig_rx =-904;
25521: waveform_sig_rx =-704;
25522: waveform_sig_rx =-761;
25523: waveform_sig_rx =-939;
25524: waveform_sig_rx =-756;
25525: waveform_sig_rx =-654;
25526: waveform_sig_rx =-871;
25527: waveform_sig_rx =-860;
25528: waveform_sig_rx =-601;
25529: waveform_sig_rx =-779;
25530: waveform_sig_rx =-941;
25531: waveform_sig_rx =-523;
25532: waveform_sig_rx =-798;
25533: waveform_sig_rx =-864;
25534: waveform_sig_rx =-616;
25535: waveform_sig_rx =-683;
25536: waveform_sig_rx =-801;
25537: waveform_sig_rx =-741;
25538: waveform_sig_rx =-560;
25539: waveform_sig_rx =-761;
25540: waveform_sig_rx =-826;
25541: waveform_sig_rx =-476;
25542: waveform_sig_rx =-744;
25543: waveform_sig_rx =-773;
25544: waveform_sig_rx =-573;
25545: waveform_sig_rx =-775;
25546: waveform_sig_rx =-596;
25547: waveform_sig_rx =-708;
25548: waveform_sig_rx =-575;
25549: waveform_sig_rx =-859;
25550: waveform_sig_rx =-423;
25551: waveform_sig_rx =-754;
25552: waveform_sig_rx =-764;
25553: waveform_sig_rx =-370;
25554: waveform_sig_rx =-814;
25555: waveform_sig_rx =-652;
25556: waveform_sig_rx =-422;
25557: waveform_sig_rx =-748;
25558: waveform_sig_rx =-648;
25559: waveform_sig_rx =-460;
25560: waveform_sig_rx =-635;
25561: waveform_sig_rx =-656;
25562: waveform_sig_rx =-496;
25563: waveform_sig_rx =-455;
25564: waveform_sig_rx =-761;
25565: waveform_sig_rx =-465;
25566: waveform_sig_rx =-407;
25567: waveform_sig_rx =-691;
25568: waveform_sig_rx =-550;
25569: waveform_sig_rx =-373;
25570: waveform_sig_rx =-574;
25571: waveform_sig_rx =-634;
25572: waveform_sig_rx =-323;
25573: waveform_sig_rx =-532;
25574: waveform_sig_rx =-608;
25575: waveform_sig_rx =-397;
25576: waveform_sig_rx =-404;
25577: waveform_sig_rx =-573;
25578: waveform_sig_rx =-495;
25579: waveform_sig_rx =-276;
25580: waveform_sig_rx =-534;
25581: waveform_sig_rx =-572;
25582: waveform_sig_rx =-192;
25583: waveform_sig_rx =-552;
25584: waveform_sig_rx =-492;
25585: waveform_sig_rx =-309;
25586: waveform_sig_rx =-569;
25587: waveform_sig_rx =-287;
25588: waveform_sig_rx =-449;
25589: waveform_sig_rx =-355;
25590: waveform_sig_rx =-540;
25591: waveform_sig_rx =-199;
25592: waveform_sig_rx =-483;
25593: waveform_sig_rx =-440;
25594: waveform_sig_rx =-154;
25595: waveform_sig_rx =-493;
25596: waveform_sig_rx =-384;
25597: waveform_sig_rx =-158;
25598: waveform_sig_rx =-431;
25599: waveform_sig_rx =-426;
25600: waveform_sig_rx =-142;
25601: waveform_sig_rx =-365;
25602: waveform_sig_rx =-438;
25603: waveform_sig_rx =-157;
25604: waveform_sig_rx =-214;
25605: waveform_sig_rx =-523;
25606: waveform_sig_rx =-142;
25607: waveform_sig_rx =-180;
25608: waveform_sig_rx =-408;
25609: waveform_sig_rx =-249;
25610: waveform_sig_rx =-148;
25611: waveform_sig_rx =-304;
25612: waveform_sig_rx =-326;
25613: waveform_sig_rx =-86;
25614: waveform_sig_rx =-221;
25615: waveform_sig_rx =-332;
25616: waveform_sig_rx =-144;
25617: waveform_sig_rx =-71;
25618: waveform_sig_rx =-343;
25619: waveform_sig_rx =-207;
25620: waveform_sig_rx =24;
25621: waveform_sig_rx =-335;
25622: waveform_sig_rx =-221;
25623: waveform_sig_rx =68;
25624: waveform_sig_rx =-307;
25625: waveform_sig_rx =-117;
25626: waveform_sig_rx =-89;
25627: waveform_sig_rx =-252;
25628: waveform_sig_rx =34;
25629: waveform_sig_rx =-223;
25630: waveform_sig_rx =-16;
25631: waveform_sig_rx =-243;
25632: waveform_sig_rx =63;
25633: waveform_sig_rx =-150;
25634: waveform_sig_rx =-178;
25635: waveform_sig_rx =142;
25636: waveform_sig_rx =-183;
25637: waveform_sig_rx =-130;
25638: waveform_sig_rx =165;
25639: waveform_sig_rx =-149;
25640: waveform_sig_rx =-156;
25641: waveform_sig_rx =183;
25642: waveform_sig_rx =-90;
25643: waveform_sig_rx =-145;
25644: waveform_sig_rx =166;
25645: waveform_sig_rx =37;
25646: waveform_sig_rx =-228;
25647: waveform_sig_rx =175;
25648: waveform_sig_rx =46;
25649: waveform_sig_rx =-81;
25650: waveform_sig_rx =57;
25651: waveform_sig_rx =129;
25652: waveform_sig_rx =27;
25653: waveform_sig_rx =-75;
25654: waveform_sig_rx =214;
25655: waveform_sig_rx =97;
25656: waveform_sig_rx =-101;
25657: waveform_sig_rx =198;
25658: waveform_sig_rx =214;
25659: waveform_sig_rx =-110;
25660: waveform_sig_rx =169;
25661: waveform_sig_rx =269;
25662: waveform_sig_rx =-53;
25663: waveform_sig_rx =132;
25664: waveform_sig_rx =292;
25665: waveform_sig_rx =31;
25666: waveform_sig_rx =168;
25667: waveform_sig_rx =161;
25668: waveform_sig_rx =137;
25669: waveform_sig_rx =258;
25670: waveform_sig_rx =84;
25671: waveform_sig_rx =307;
25672: waveform_sig_rx =7;
25673: waveform_sig_rx =402;
25674: waveform_sig_rx =126;
25675: waveform_sig_rx =99;
25676: waveform_sig_rx =436;
25677: waveform_sig_rx =79;
25678: waveform_sig_rx =154;
25679: waveform_sig_rx =474;
25680: waveform_sig_rx =112;
25681: waveform_sig_rx =156;
25682: waveform_sig_rx =538;
25683: waveform_sig_rx =128;
25684: waveform_sig_rx =192;
25685: waveform_sig_rx =479;
25686: waveform_sig_rx =248;
25687: waveform_sig_rx =160;
25688: waveform_sig_rx =442;
25689: waveform_sig_rx =341;
25690: waveform_sig_rx =277;
25691: waveform_sig_rx =277;
25692: waveform_sig_rx =475;
25693: waveform_sig_rx =296;
25694: waveform_sig_rx =199;
25695: waveform_sig_rx =565;
25696: waveform_sig_rx =311;
25697: waveform_sig_rx =216;
25698: waveform_sig_rx =523;
25699: waveform_sig_rx =420;
25700: waveform_sig_rx =199;
25701: waveform_sig_rx =464;
25702: waveform_sig_rx =503;
25703: waveform_sig_rx =257;
25704: waveform_sig_rx =407;
25705: waveform_sig_rx =561;
25706: waveform_sig_rx =353;
25707: waveform_sig_rx =426;
25708: waveform_sig_rx =425;
25709: waveform_sig_rx =455;
25710: waveform_sig_rx =475;
25711: waveform_sig_rx =414;
25712: waveform_sig_rx =563;
25713: waveform_sig_rx =256;
25714: waveform_sig_rx =716;
25715: waveform_sig_rx =367;
25716: waveform_sig_rx =369;
25717: waveform_sig_rx =760;
25718: waveform_sig_rx =296;
25719: waveform_sig_rx =481;
25720: waveform_sig_rx =777;
25721: waveform_sig_rx =325;
25722: waveform_sig_rx =477;
25723: waveform_sig_rx =768;
25724: waveform_sig_rx =365;
25725: waveform_sig_rx =498;
25726: waveform_sig_rx =669;
25727: waveform_sig_rx =549;
25728: waveform_sig_rx =434;
25729: waveform_sig_rx =674;
25730: waveform_sig_rx =641;
25731: waveform_sig_rx =488;
25732: waveform_sig_rx =532;
25733: waveform_sig_rx =799;
25734: waveform_sig_rx =486;
25735: waveform_sig_rx =524;
25736: waveform_sig_rx =842;
25737: waveform_sig_rx =539;
25738: waveform_sig_rx =529;
25739: waveform_sig_rx =777;
25740: waveform_sig_rx =661;
25741: waveform_sig_rx =501;
25742: waveform_sig_rx =725;
25743: waveform_sig_rx =753;
25744: waveform_sig_rx =557;
25745: waveform_sig_rx =617;
25746: waveform_sig_rx =840;
25747: waveform_sig_rx =609;
25748: waveform_sig_rx =642;
25749: waveform_sig_rx =745;
25750: waveform_sig_rx =672;
25751: waveform_sig_rx =716;
25752: waveform_sig_rx =723;
25753: waveform_sig_rx =725;
25754: waveform_sig_rx =549;
25755: waveform_sig_rx =989;
25756: waveform_sig_rx =525;
25757: waveform_sig_rx =724;
25758: waveform_sig_rx =945;
25759: waveform_sig_rx =518;
25760: waveform_sig_rx =778;
25761: waveform_sig_rx =952;
25762: waveform_sig_rx =568;
25763: waveform_sig_rx =746;
25764: waveform_sig_rx =975;
25765: waveform_sig_rx =647;
25766: waveform_sig_rx =774;
25767: waveform_sig_rx =883;
25768: waveform_sig_rx =812;
25769: waveform_sig_rx =638;
25770: waveform_sig_rx =912;
25771: waveform_sig_rx =904;
25772: waveform_sig_rx =676;
25773: waveform_sig_rx =799;
25774: waveform_sig_rx =1030;
25775: waveform_sig_rx =676;
25776: waveform_sig_rx =808;
25777: waveform_sig_rx =1023;
25778: waveform_sig_rx =767;
25779: waveform_sig_rx =804;
25780: waveform_sig_rx =952;
25781: waveform_sig_rx =926;
25782: waveform_sig_rx =723;
25783: waveform_sig_rx =889;
25784: waveform_sig_rx =1018;
25785: waveform_sig_rx =742;
25786: waveform_sig_rx =842;
25787: waveform_sig_rx =1113;
25788: waveform_sig_rx =761;
25789: waveform_sig_rx =886;
25790: waveform_sig_rx =985;
25791: waveform_sig_rx =842;
25792: waveform_sig_rx =964;
25793: waveform_sig_rx =928;
25794: waveform_sig_rx =904;
25795: waveform_sig_rx =802;
25796: waveform_sig_rx =1123;
25797: waveform_sig_rx =724;
25798: waveform_sig_rx =970;
25799: waveform_sig_rx =1080;
25800: waveform_sig_rx =734;
25801: waveform_sig_rx =961;
25802: waveform_sig_rx =1120;
25803: waveform_sig_rx =775;
25804: waveform_sig_rx =925;
25805: waveform_sig_rx =1141;
25806: waveform_sig_rx =842;
25807: waveform_sig_rx =933;
25808: waveform_sig_rx =1077;
25809: waveform_sig_rx =1016;
25810: waveform_sig_rx =745;
25811: waveform_sig_rx =1136;
25812: waveform_sig_rx =1069;
25813: waveform_sig_rx =785;
25814: waveform_sig_rx =1081;
25815: waveform_sig_rx =1123;
25816: waveform_sig_rx =855;
25817: waveform_sig_rx =1045;
25818: waveform_sig_rx =1106;
25819: waveform_sig_rx =1012;
25820: waveform_sig_rx =918;
25821: waveform_sig_rx =1108;
25822: waveform_sig_rx =1155;
25823: waveform_sig_rx =812;
25824: waveform_sig_rx =1148;
25825: waveform_sig_rx =1176;
25826: waveform_sig_rx =850;
25827: waveform_sig_rx =1080;
25828: waveform_sig_rx =1206;
25829: waveform_sig_rx =905;
25830: waveform_sig_rx =1087;
25831: waveform_sig_rx =1077;
25832: waveform_sig_rx =1015;
25833: waveform_sig_rx =1115;
25834: waveform_sig_rx =1054;
25835: waveform_sig_rx =1045;
25836: waveform_sig_rx =996;
25837: waveform_sig_rx =1253;
25838: waveform_sig_rx =886;
25839: waveform_sig_rx =1127;
25840: waveform_sig_rx =1174;
25841: waveform_sig_rx =944;
25842: waveform_sig_rx =1094;
25843: waveform_sig_rx =1238;
25844: waveform_sig_rx =953;
25845: waveform_sig_rx =996;
25846: waveform_sig_rx =1342;
25847: waveform_sig_rx =931;
25848: waveform_sig_rx =1029;
25849: waveform_sig_rx =1296;
25850: waveform_sig_rx =1031;
25851: waveform_sig_rx =932;
25852: waveform_sig_rx =1312;
25853: waveform_sig_rx =1091;
25854: waveform_sig_rx =1011;
25855: waveform_sig_rx =1153;
25856: waveform_sig_rx =1216;
25857: waveform_sig_rx =1021;
25858: waveform_sig_rx =1080;
25859: waveform_sig_rx =1265;
25860: waveform_sig_rx =1110;
25861: waveform_sig_rx =978;
25862: waveform_sig_rx =1265;
25863: waveform_sig_rx =1194;
25864: waveform_sig_rx =893;
25865: waveform_sig_rx =1272;
25866: waveform_sig_rx =1227;
25867: waveform_sig_rx =942;
25868: waveform_sig_rx =1202;
25869: waveform_sig_rx =1277;
25870: waveform_sig_rx =984;
25871: waveform_sig_rx =1219;
25872: waveform_sig_rx =1084;
25873: waveform_sig_rx =1127;
25874: waveform_sig_rx =1205;
25875: waveform_sig_rx =1101;
25876: waveform_sig_rx =1178;
25877: waveform_sig_rx =1048;
25878: waveform_sig_rx =1313;
25879: waveform_sig_rx =999;
25880: waveform_sig_rx =1149;
25881: waveform_sig_rx =1303;
25882: waveform_sig_rx =1012;
25883: waveform_sig_rx =1107;
25884: waveform_sig_rx =1398;
25885: waveform_sig_rx =932;
25886: waveform_sig_rx =1114;
25887: waveform_sig_rx =1440;
25888: waveform_sig_rx =900;
25889: waveform_sig_rx =1189;
25890: waveform_sig_rx =1314;
25891: waveform_sig_rx =1048;
25892: waveform_sig_rx =1066;
25893: waveform_sig_rx =1307;
25894: waveform_sig_rx =1144;
25895: waveform_sig_rx =1067;
25896: waveform_sig_rx =1163;
25897: waveform_sig_rx =1306;
25898: waveform_sig_rx =1024;
25899: waveform_sig_rx =1117;
25900: waveform_sig_rx =1324;
25901: waveform_sig_rx =1069;
25902: waveform_sig_rx =1024;
25903: waveform_sig_rx =1318;
25904: waveform_sig_rx =1181;
25905: waveform_sig_rx =939;
25906: waveform_sig_rx =1326;
25907: waveform_sig_rx =1191;
25908: waveform_sig_rx =979;
25909: waveform_sig_rx =1237;
25910: waveform_sig_rx =1221;
25911: waveform_sig_rx =1037;
25912: waveform_sig_rx =1196;
25913: waveform_sig_rx =1069;
25914: waveform_sig_rx =1226;
25915: waveform_sig_rx =1111;
25916: waveform_sig_rx =1156;
25917: waveform_sig_rx =1180;
25918: waveform_sig_rx =970;
25919: waveform_sig_rx =1385;
25920: waveform_sig_rx =929;
25921: waveform_sig_rx =1117;
25922: waveform_sig_rx =1353;
25923: waveform_sig_rx =879;
25924: waveform_sig_rx =1199;
25925: waveform_sig_rx =1338;
25926: waveform_sig_rx =860;
25927: waveform_sig_rx =1188;
25928: waveform_sig_rx =1325;
25929: waveform_sig_rx =915;
25930: waveform_sig_rx =1179;
25931: waveform_sig_rx =1231;
25932: waveform_sig_rx =1064;
25933: waveform_sig_rx =1006;
25934: waveform_sig_rx =1268;
25935: waveform_sig_rx =1124;
25936: waveform_sig_rx =1032;
25937: waveform_sig_rx =1118;
25938: waveform_sig_rx =1270;
25939: waveform_sig_rx =972;
25940: waveform_sig_rx =1077;
25941: waveform_sig_rx =1315;
25942: waveform_sig_rx =985;
25943: waveform_sig_rx =994;
25944: waveform_sig_rx =1297;
25945: waveform_sig_rx =1039;
25946: waveform_sig_rx =983;
25947: waveform_sig_rx =1230;
25948: waveform_sig_rx =1093;
25949: waveform_sig_rx =1020;
25950: waveform_sig_rx =1072;
25951: waveform_sig_rx =1224;
25952: waveform_sig_rx =974;
25953: waveform_sig_rx =1079;
25954: waveform_sig_rx =1077;
25955: waveform_sig_rx =1092;
25956: waveform_sig_rx =1035;
25957: waveform_sig_rx =1149;
25958: waveform_sig_rx =1040;
25959: waveform_sig_rx =976;
25960: waveform_sig_rx =1334;
25961: waveform_sig_rx =791;
25962: waveform_sig_rx =1148;
25963: waveform_sig_rx =1197;
25964: waveform_sig_rx =780;
25965: waveform_sig_rx =1184;
25966: waveform_sig_rx =1197;
25967: waveform_sig_rx =800;
25968: waveform_sig_rx =1152;
25969: waveform_sig_rx =1190;
25970: waveform_sig_rx =859;
25971: waveform_sig_rx =1086;
25972: waveform_sig_rx =1114;
25973: waveform_sig_rx =990;
25974: waveform_sig_rx =859;
25975: waveform_sig_rx =1151;
25976: waveform_sig_rx =1015;
25977: waveform_sig_rx =868;
25978: waveform_sig_rx =1018;
25979: waveform_sig_rx =1157;
25980: waveform_sig_rx =790;
25981: waveform_sig_rx =1010;
25982: waveform_sig_rx =1163;
25983: waveform_sig_rx =825;
25984: waveform_sig_rx =934;
25985: waveform_sig_rx =1106;
25986: waveform_sig_rx =939;
25987: waveform_sig_rx =867;
25988: waveform_sig_rx =1038;
25989: waveform_sig_rx =1053;
25990: waveform_sig_rx =822;
25991: waveform_sig_rx =963;
25992: waveform_sig_rx =1161;
25993: waveform_sig_rx =754;
25994: waveform_sig_rx =1036;
25995: waveform_sig_rx =943;
25996: waveform_sig_rx =919;
25997: waveform_sig_rx =981;
25998: waveform_sig_rx =976;
25999: waveform_sig_rx =869;
26000: waveform_sig_rx =893;
26001: waveform_sig_rx =1104;
26002: waveform_sig_rx =659;
26003: waveform_sig_rx =1030;
26004: waveform_sig_rx =984;
26005: waveform_sig_rx =668;
26006: waveform_sig_rx =1022;
26007: waveform_sig_rx =977;
26008: waveform_sig_rx =668;
26009: waveform_sig_rx =951;
26010: waveform_sig_rx =987;
26011: waveform_sig_rx =724;
26012: waveform_sig_rx =862;
26013: waveform_sig_rx =962;
26014: waveform_sig_rx =809;
26015: waveform_sig_rx =652;
26016: waveform_sig_rx =1051;
26017: waveform_sig_rx =793;
26018: waveform_sig_rx =690;
26019: waveform_sig_rx =922;
26020: waveform_sig_rx =914;
26021: waveform_sig_rx =659;
26022: waveform_sig_rx =873;
26023: waveform_sig_rx =910;
26024: waveform_sig_rx =696;
26025: waveform_sig_rx =741;
26026: waveform_sig_rx =907;
26027: waveform_sig_rx =788;
26028: waveform_sig_rx =632;
26029: waveform_sig_rx =894;
26030: waveform_sig_rx =855;
26031: waveform_sig_rx =578;
26032: waveform_sig_rx =846;
26033: waveform_sig_rx =910;
26034: waveform_sig_rx =522;
26035: waveform_sig_rx =904;
26036: waveform_sig_rx =656;
26037: waveform_sig_rx =757;
26038: waveform_sig_rx =749;
26039: waveform_sig_rx =701;
26040: waveform_sig_rx =670;
26041: waveform_sig_rx =677;
26042: waveform_sig_rx =849;
26043: waveform_sig_rx =491;
26044: waveform_sig_rx =790;
26045: waveform_sig_rx =767;
26046: waveform_sig_rx =498;
26047: waveform_sig_rx =783;
26048: waveform_sig_rx =778;
26049: waveform_sig_rx =481;
26050: waveform_sig_rx =701;
26051: waveform_sig_rx =808;
26052: waveform_sig_rx =487;
26053: waveform_sig_rx =644;
26054: waveform_sig_rx =811;
26055: waveform_sig_rx =525;
26056: waveform_sig_rx =489;
26057: waveform_sig_rx =849;
26058: waveform_sig_rx =514;
26059: waveform_sig_rx =545;
26060: waveform_sig_rx =660;
26061: waveform_sig_rx =673;
26062: waveform_sig_rx =469;
26063: waveform_sig_rx =600;
26064: waveform_sig_rx =691;
26065: waveform_sig_rx =473;
26066: waveform_sig_rx =475;
26067: waveform_sig_rx =705;
26068: waveform_sig_rx =542;
26069: waveform_sig_rx =355;
26070: waveform_sig_rx =721;
26071: waveform_sig_rx =558;
26072: waveform_sig_rx =306;
26073: waveform_sig_rx =647;
26074: waveform_sig_rx =572;
26075: waveform_sig_rx =315;
26076: waveform_sig_rx =630;
26077: waveform_sig_rx =327;
26078: waveform_sig_rx =574;
26079: waveform_sig_rx =438;
26080: waveform_sig_rx =472;
26081: waveform_sig_rx =464;
26082: waveform_sig_rx =367;
26083: waveform_sig_rx =625;
26084: waveform_sig_rx =221;
26085: waveform_sig_rx =515;
26086: waveform_sig_rx =538;
26087: waveform_sig_rx =181;
26088: waveform_sig_rx =538;
26089: waveform_sig_rx =519;
26090: waveform_sig_rx =177;
26091: waveform_sig_rx =469;
26092: waveform_sig_rx =545;
26093: waveform_sig_rx =180;
26094: waveform_sig_rx =383;
26095: waveform_sig_rx =539;
26096: waveform_sig_rx =196;
26097: waveform_sig_rx =275;
26098: waveform_sig_rx =552;
26099: waveform_sig_rx =214;
26100: waveform_sig_rx =322;
26101: waveform_sig_rx =340;
26102: waveform_sig_rx =432;
26103: waveform_sig_rx =185;
26104: waveform_sig_rx =273;
26105: waveform_sig_rx =475;
26106: waveform_sig_rx =134;
26107: waveform_sig_rx =206;
26108: waveform_sig_rx =468;
26109: waveform_sig_rx =143;
26110: waveform_sig_rx =132;
26111: waveform_sig_rx =401;
26112: waveform_sig_rx =203;
26113: waveform_sig_rx =101;
26114: waveform_sig_rx =304;
26115: waveform_sig_rx =295;
26116: waveform_sig_rx =79;
26117: waveform_sig_rx =286;
26118: waveform_sig_rx =94;
26119: waveform_sig_rx =294;
26120: waveform_sig_rx =115;
26121: waveform_sig_rx =242;
26122: waveform_sig_rx =109;
26123: waveform_sig_rx =95;
26124: waveform_sig_rx =352;
26125: waveform_sig_rx =-114;
26126: waveform_sig_rx =255;
26127: waveform_sig_rx =236;
26128: waveform_sig_rx =-143;
26129: waveform_sig_rx =274;
26130: waveform_sig_rx =211;
26131: waveform_sig_rx =-161;
26132: waveform_sig_rx =238;
26133: waveform_sig_rx =207;
26134: waveform_sig_rx =-161;
26135: waveform_sig_rx =171;
26136: waveform_sig_rx =178;
26137: waveform_sig_rx =-99;
26138: waveform_sig_rx =8;
26139: waveform_sig_rx =172;
26140: waveform_sig_rx =-21;
26141: waveform_sig_rx =-37;
26142: waveform_sig_rx =-2;
26143: waveform_sig_rx =192;
26144: waveform_sig_rx =-219;
26145: waveform_sig_rx =30;
26146: waveform_sig_rx =181;
26147: waveform_sig_rx =-241;
26148: waveform_sig_rx =-9;
26149: waveform_sig_rx =115;
26150: waveform_sig_rx =-152;
26151: waveform_sig_rx =-106;
26152: waveform_sig_rx =65;
26153: waveform_sig_rx =-61;
26154: waveform_sig_rx =-207;
26155: waveform_sig_rx =-12;
26156: waveform_sig_rx =15;
26157: waveform_sig_rx =-274;
26158: waveform_sig_rx =-13;
26159: waveform_sig_rx =-202;
26160: waveform_sig_rx =-46;
26161: waveform_sig_rx =-191;
26162: waveform_sig_rx =-49;
26163: waveform_sig_rx =-236;
26164: waveform_sig_rx =-181;
26165: waveform_sig_rx =39;
26166: waveform_sig_rx =-439;
26167: waveform_sig_rx =-20;
26168: waveform_sig_rx =-79;
26169: waveform_sig_rx =-476;
26170: waveform_sig_rx =31;
26171: waveform_sig_rx =-161;
26172: waveform_sig_rx =-471;
26173: waveform_sig_rx =-35;
26174: waveform_sig_rx =-214;
26175: waveform_sig_rx =-393;
26176: waveform_sig_rx =-183;
26177: waveform_sig_rx =-178;
26178: waveform_sig_rx =-319;
26179: waveform_sig_rx =-387;
26180: waveform_sig_rx =-101;
26181: waveform_sig_rx =-327;
26182: waveform_sig_rx =-408;
26183: waveform_sig_rx =-202;
26184: waveform_sig_rx =-186;
26185: waveform_sig_rx =-520;
26186: waveform_sig_rx =-203;
26187: waveform_sig_rx =-210;
26188: waveform_sig_rx =-499;
26189: waveform_sig_rx =-323;
26190: waveform_sig_rx =-203;
26191: waveform_sig_rx =-444;
26192: waveform_sig_rx =-444;
26193: waveform_sig_rx =-228;
26194: waveform_sig_rx =-380;
26195: waveform_sig_rx =-526;
26196: waveform_sig_rx =-332;
26197: waveform_sig_rx =-265;
26198: waveform_sig_rx =-571;
26199: waveform_sig_rx =-309;
26200: waveform_sig_rx =-445;
26201: waveform_sig_rx =-385;
26202: waveform_sig_rx =-458;
26203: waveform_sig_rx =-319;
26204: waveform_sig_rx =-588;
26205: waveform_sig_rx =-369;
26206: waveform_sig_rx =-332;
26207: waveform_sig_rx =-736;
26208: waveform_sig_rx =-235;
26209: waveform_sig_rx =-493;
26210: waveform_sig_rx =-671;
26211: waveform_sig_rx =-292;
26212: waveform_sig_rx =-498;
26213: waveform_sig_rx =-680;
26214: waveform_sig_rx =-386;
26215: waveform_sig_rx =-452;
26216: waveform_sig_rx =-669;
26217: waveform_sig_rx =-489;
26218: waveform_sig_rx =-418;
26219: waveform_sig_rx =-656;
26220: waveform_sig_rx =-641;
26221: waveform_sig_rx =-351;
26222: waveform_sig_rx =-636;
26223: waveform_sig_rx =-676;
26224: waveform_sig_rx =-457;
26225: waveform_sig_rx =-502;
26226: waveform_sig_rx =-792;
26227: waveform_sig_rx =-459;
26228: waveform_sig_rx =-537;
26229: waveform_sig_rx =-749;
26230: waveform_sig_rx =-598;
26231: waveform_sig_rx =-511;
26232: waveform_sig_rx =-672;
26233: waveform_sig_rx =-764;
26234: waveform_sig_rx =-491;
26235: waveform_sig_rx =-615;
26236: waveform_sig_rx =-828;
26237: waveform_sig_rx =-528;
26238: waveform_sig_rx =-569;
26239: waveform_sig_rx =-877;
26240: waveform_sig_rx =-533;
26241: waveform_sig_rx =-775;
26242: waveform_sig_rx =-647;
26243: waveform_sig_rx =-680;
26244: waveform_sig_rx =-652;
26245: waveform_sig_rx =-841;
26246: waveform_sig_rx =-627;
26247: waveform_sig_rx =-691;
26248: waveform_sig_rx =-925;
26249: waveform_sig_rx =-542;
26250: waveform_sig_rx =-789;
26251: waveform_sig_rx =-873;
26252: waveform_sig_rx =-609;
26253: waveform_sig_rx =-713;
26254: waveform_sig_rx =-950;
26255: waveform_sig_rx =-673;
26256: waveform_sig_rx =-662;
26257: waveform_sig_rx =-971;
26258: waveform_sig_rx =-716;
26259: waveform_sig_rx =-665;
26260: waveform_sig_rx =-949;
26261: waveform_sig_rx =-879;
26262: waveform_sig_rx =-615;
26263: waveform_sig_rx =-920;
26264: waveform_sig_rx =-924;
26265: waveform_sig_rx =-696;
26266: waveform_sig_rx =-806;
26267: waveform_sig_rx =-991;
26268: waveform_sig_rx =-722;
26269: waveform_sig_rx =-786;
26270: waveform_sig_rx =-929;
26271: waveform_sig_rx =-911;
26272: waveform_sig_rx =-698;
26273: waveform_sig_rx =-904;
26274: waveform_sig_rx =-1050;
26275: waveform_sig_rx =-642;
26276: waveform_sig_rx =-942;
26277: waveform_sig_rx =-1054;
26278: waveform_sig_rx =-713;
26279: waveform_sig_rx =-902;
26280: waveform_sig_rx =-1038;
26281: waveform_sig_rx =-794;
26282: waveform_sig_rx =-1049;
26283: waveform_sig_rx =-820;
26284: waveform_sig_rx =-993;
26285: waveform_sig_rx =-870;
26286: waveform_sig_rx =-1037;
26287: waveform_sig_rx =-852;
26288: waveform_sig_rx =-888;
26289: waveform_sig_rx =-1119;
26290: waveform_sig_rx =-793;
26291: waveform_sig_rx =-975;
26292: waveform_sig_rx =-1110;
26293: waveform_sig_rx =-837;
26294: waveform_sig_rx =-893;
26295: waveform_sig_rx =-1205;
26296: waveform_sig_rx =-849;
26297: waveform_sig_rx =-872;
26298: waveform_sig_rx =-1245;
26299: waveform_sig_rx =-862;
26300: waveform_sig_rx =-858;
26301: waveform_sig_rx =-1186;
26302: waveform_sig_rx =-980;
26303: waveform_sig_rx =-861;
26304: waveform_sig_rx =-1138;
26305: waveform_sig_rx =-1041;
26306: waveform_sig_rx =-950;
26307: waveform_sig_rx =-962;
26308: waveform_sig_rx =-1173;
26309: waveform_sig_rx =-948;
26310: waveform_sig_rx =-934;
26311: waveform_sig_rx =-1176;
26312: waveform_sig_rx =-1080;
26313: waveform_sig_rx =-849;
26314: waveform_sig_rx =-1169;
26315: waveform_sig_rx =-1154;
26316: waveform_sig_rx =-825;
26317: waveform_sig_rx =-1153;
26318: waveform_sig_rx =-1157;
26319: waveform_sig_rx =-909;
26320: waveform_sig_rx =-1054;
26321: waveform_sig_rx =-1150;
26322: waveform_sig_rx =-978;
26323: waveform_sig_rx =-1196;
26324: waveform_sig_rx =-974;
26325: waveform_sig_rx =-1161;
26326: waveform_sig_rx =-1017;
26327: waveform_sig_rx =-1216;
26328: waveform_sig_rx =-1051;
26329: waveform_sig_rx =-1029;
26330: waveform_sig_rx =-1284;
26331: waveform_sig_rx =-982;
26332: waveform_sig_rx =-1073;
26333: waveform_sig_rx =-1299;
26334: waveform_sig_rx =-941;
26335: waveform_sig_rx =-1037;
26336: waveform_sig_rx =-1404;
26337: waveform_sig_rx =-880;
26338: waveform_sig_rx =-1076;
26339: waveform_sig_rx =-1351;
26340: waveform_sig_rx =-932;
26341: waveform_sig_rx =-1081;
26342: waveform_sig_rx =-1256;
26343: waveform_sig_rx =-1100;
26344: waveform_sig_rx =-1013;
26345: waveform_sig_rx =-1188;
26346: waveform_sig_rx =-1215;
26347: waveform_sig_rx =-1058;
26348: waveform_sig_rx =-1060;
26349: waveform_sig_rx =-1322;
26350: waveform_sig_rx =-1028;
26351: waveform_sig_rx =-1044;
26352: waveform_sig_rx =-1309;
26353: waveform_sig_rx =-1128;
26354: waveform_sig_rx =-973;
26355: waveform_sig_rx =-1304;
26356: waveform_sig_rx =-1190;
26357: waveform_sig_rx =-973;
26358: waveform_sig_rx =-1256;
26359: waveform_sig_rx =-1211;
26360: waveform_sig_rx =-1047;
26361: waveform_sig_rx =-1129;
26362: waveform_sig_rx =-1231;
26363: waveform_sig_rx =-1105;
26364: waveform_sig_rx =-1212;
26365: waveform_sig_rx =-1049;
26366: waveform_sig_rx =-1265;
26367: waveform_sig_rx =-1018;
26368: waveform_sig_rx =-1325;
26369: waveform_sig_rx =-1077;
26370: waveform_sig_rx =-1059;
26371: waveform_sig_rx =-1400;
26372: waveform_sig_rx =-943;
26373: waveform_sig_rx =-1174;
26374: waveform_sig_rx =-1377;
26375: waveform_sig_rx =-908;
26376: waveform_sig_rx =-1180;
26377: waveform_sig_rx =-1370;
26378: waveform_sig_rx =-935;
26379: waveform_sig_rx =-1211;
26380: waveform_sig_rx =-1310;
26381: waveform_sig_rx =-1025;
26382: waveform_sig_rx =-1131;
26383: waveform_sig_rx =-1278;
26384: waveform_sig_rx =-1198;
26385: waveform_sig_rx =-1035;
26386: waveform_sig_rx =-1231;
26387: waveform_sig_rx =-1267;
26388: waveform_sig_rx =-1048;
26389: waveform_sig_rx =-1129;
26390: waveform_sig_rx =-1356;
26391: waveform_sig_rx =-1005;
26392: waveform_sig_rx =-1091;
26393: waveform_sig_rx =-1345;
26394: waveform_sig_rx =-1090;
26395: waveform_sig_rx =-1027;
26396: waveform_sig_rx =-1315;
26397: waveform_sig_rx =-1148;
26398: waveform_sig_rx =-1036;
26399: waveform_sig_rx =-1222;
26400: waveform_sig_rx =-1230;
26401: waveform_sig_rx =-1094;
26402: waveform_sig_rx =-1074;
26403: waveform_sig_rx =-1288;
26404: waveform_sig_rx =-1080;
26405: waveform_sig_rx =-1187;
26406: waveform_sig_rx =-1130;
26407: waveform_sig_rx =-1187;
26408: waveform_sig_rx =-1033;
26409: waveform_sig_rx =-1341;
26410: waveform_sig_rx =-962;
26411: waveform_sig_rx =-1145;
26412: waveform_sig_rx =-1343;
26413: waveform_sig_rx =-882;
26414: waveform_sig_rx =-1237;
26415: waveform_sig_rx =-1273;
26416: waveform_sig_rx =-915;
26417: waveform_sig_rx =-1179;
26418: waveform_sig_rx =-1296;
26419: waveform_sig_rx =-923;
26420: waveform_sig_rx =-1152;
26421: waveform_sig_rx =-1257;
26422: waveform_sig_rx =-1009;
26423: waveform_sig_rx =-1080;
26424: waveform_sig_rx =-1228;
26425: waveform_sig_rx =-1141;
26426: waveform_sig_rx =-962;
26427: waveform_sig_rx =-1189;
26428: waveform_sig_rx =-1234;
26429: waveform_sig_rx =-930;
26430: waveform_sig_rx =-1104;
26431: waveform_sig_rx =-1303;
26432: waveform_sig_rx =-899;
26433: waveform_sig_rx =-1127;
26434: waveform_sig_rx =-1230;
26435: waveform_sig_rx =-1036;
26436: waveform_sig_rx =-1033;
26437: waveform_sig_rx =-1174;
26438: waveform_sig_rx =-1157;
26439: waveform_sig_rx =-922;
26440: waveform_sig_rx =-1113;
26441: waveform_sig_rx =-1229;
26442: waveform_sig_rx =-902;
26443: waveform_sig_rx =-1042;
26444: waveform_sig_rx =-1225;
26445: waveform_sig_rx =-937;
26446: waveform_sig_rx =-1166;
26447: waveform_sig_rx =-1006;
26448: waveform_sig_rx =-1071;
26449: waveform_sig_rx =-994;
26450: waveform_sig_rx =-1237;
26451: waveform_sig_rx =-876;
26452: waveform_sig_rx =-1101;
26453: waveform_sig_rx =-1179;
26454: waveform_sig_rx =-814;
26455: waveform_sig_rx =-1145;
26456: waveform_sig_rx =-1116;
26457: waveform_sig_rx =-830;
26458: waveform_sig_rx =-1094;
26459: waveform_sig_rx =-1162;
26460: waveform_sig_rx =-853;
26461: waveform_sig_rx =-1025;
26462: waveform_sig_rx =-1148;
26463: waveform_sig_rx =-933;
26464: waveform_sig_rx =-909;
26465: waveform_sig_rx =-1184;
26466: waveform_sig_rx =-1004;
26467: waveform_sig_rx =-813;
26468: waveform_sig_rx =-1155;
26469: waveform_sig_rx =-1038;
26470: waveform_sig_rx =-828;
26471: waveform_sig_rx =-1042;
26472: waveform_sig_rx =-1084;
26473: waveform_sig_rx =-838;
26474: waveform_sig_rx =-977;
26475: waveform_sig_rx =-1059;
26476: waveform_sig_rx =-947;
26477: waveform_sig_rx =-812;
26478: waveform_sig_rx =-1063;
26479: waveform_sig_rx =-1030;
26480: waveform_sig_rx =-734;
26481: waveform_sig_rx =-1032;
26482: waveform_sig_rx =-1068;
26483: waveform_sig_rx =-690;
26484: waveform_sig_rx =-977;
26485: waveform_sig_rx =-1022;
26486: waveform_sig_rx =-756;
26487: waveform_sig_rx =-1038;
26488: waveform_sig_rx =-773;
26489: waveform_sig_rx =-938;
26490: waveform_sig_rx =-829;
26491: waveform_sig_rx =-1012;
26492: waveform_sig_rx =-708;
26493: waveform_sig_rx =-931;
26494: waveform_sig_rx =-988;
26495: waveform_sig_rx =-693;
26496: waveform_sig_rx =-953;
26497: waveform_sig_rx =-958;
26498: waveform_sig_rx =-681;
26499: waveform_sig_rx =-872;
26500: waveform_sig_rx =-995;
26501: waveform_sig_rx =-665;
26502: waveform_sig_rx =-836;
26503: waveform_sig_rx =-1005;
26504: waveform_sig_rx =-726;
26505: waveform_sig_rx =-719;
26506: waveform_sig_rx =-1037;
26507: waveform_sig_rx =-721;
26508: waveform_sig_rx =-678;
26509: waveform_sig_rx =-954;
26510: waveform_sig_rx =-774;
26511: waveform_sig_rx =-711;
26512: waveform_sig_rx =-764;
26513: waveform_sig_rx =-888;
26514: waveform_sig_rx =-686;
26515: waveform_sig_rx =-706;
26516: waveform_sig_rx =-902;
26517: waveform_sig_rx =-702;
26518: waveform_sig_rx =-585;
26519: waveform_sig_rx =-925;
26520: waveform_sig_rx =-770;
26521: waveform_sig_rx =-523;
26522: waveform_sig_rx =-873;
26523: waveform_sig_rx =-784;
26524: waveform_sig_rx =-520;
26525: waveform_sig_rx =-796;
26526: waveform_sig_rx =-733;
26527: waveform_sig_rx =-615;
26528: waveform_sig_rx =-822;
26529: waveform_sig_rx =-528;
26530: waveform_sig_rx =-786;
26531: waveform_sig_rx =-573;
26532: waveform_sig_rx =-796;
26533: waveform_sig_rx =-535;
26534: waveform_sig_rx =-647;
26535: waveform_sig_rx =-796;
26536: waveform_sig_rx =-447;
26537: waveform_sig_rx =-686;
26538: waveform_sig_rx =-759;
26539: waveform_sig_rx =-387;
26540: waveform_sig_rx =-681;
26541: waveform_sig_rx =-781;
26542: waveform_sig_rx =-359;
26543: waveform_sig_rx =-651;
26544: waveform_sig_rx =-749;
26545: waveform_sig_rx =-436;
26546: waveform_sig_rx =-525;
26547: waveform_sig_rx =-779;
26548: waveform_sig_rx =-426;
26549: waveform_sig_rx =-482;
26550: waveform_sig_rx =-651;
26551: waveform_sig_rx =-522;
26552: waveform_sig_rx =-484;
26553: waveform_sig_rx =-459;
26554: waveform_sig_rx =-702;
26555: waveform_sig_rx =-376;
26556: waveform_sig_rx =-417;
26557: waveform_sig_rx =-723;
26558: waveform_sig_rx =-360;
26559: waveform_sig_rx =-367;
26560: waveform_sig_rx =-684;
26561: waveform_sig_rx =-418;
26562: waveform_sig_rx =-351;
26563: waveform_sig_rx =-557;
26564: waveform_sig_rx =-502;
26565: waveform_sig_rx =-307;
26566: waveform_sig_rx =-464;
26567: waveform_sig_rx =-494;
26568: waveform_sig_rx =-374;
26569: waveform_sig_rx =-504;
26570: waveform_sig_rx =-314;
26571: waveform_sig_rx =-515;
26572: waveform_sig_rx =-274;
26573: waveform_sig_rx =-558;
26574: waveform_sig_rx =-213;
26575: waveform_sig_rx =-383;
26576: waveform_sig_rx =-522;
26577: waveform_sig_rx =-129;
26578: waveform_sig_rx =-464;
26579: waveform_sig_rx =-490;
26580: waveform_sig_rx =-74;
26581: waveform_sig_rx =-465;
26582: waveform_sig_rx =-479;
26583: waveform_sig_rx =-58;
26584: waveform_sig_rx =-440;
26585: waveform_sig_rx =-407;
26586: waveform_sig_rx =-160;
26587: waveform_sig_rx =-291;
26588: waveform_sig_rx =-452;
26589: waveform_sig_rx =-195;
26590: waveform_sig_rx =-220;
26591: waveform_sig_rx =-340;
26592: waveform_sig_rx =-328;
26593: waveform_sig_rx =-138;
26594: waveform_sig_rx =-238;
26595: waveform_sig_rx =-458;
26596: waveform_sig_rx =-5;
26597: waveform_sig_rx =-246;
26598: waveform_sig_rx =-388;
26599: waveform_sig_rx =-48;
26600: waveform_sig_rx =-168;
26601: waveform_sig_rx =-315;
26602: waveform_sig_rx =-166;
26603: waveform_sig_rx =-68;
26604: waveform_sig_rx =-250;
26605: waveform_sig_rx =-264;
26606: waveform_sig_rx =4;
26607: waveform_sig_rx =-215;
26608: waveform_sig_rx =-224;
26609: waveform_sig_rx =-80;
26610: waveform_sig_rx =-214;
26611: waveform_sig_rx =-61;
26612: waveform_sig_rx =-207;
26613: waveform_sig_rx =-2;
26614: waveform_sig_rx =-301;
26615: waveform_sig_rx =112;
26616: waveform_sig_rx =-158;
26617: waveform_sig_rx =-243;
26618: waveform_sig_rx =199;
26619: waveform_sig_rx =-236;
26620: waveform_sig_rx =-153;
26621: waveform_sig_rx =230;
26622: waveform_sig_rx =-231;
26623: waveform_sig_rx =-101;
26624: waveform_sig_rx =161;
26625: waveform_sig_rx =-164;
26626: waveform_sig_rx =-58;
26627: waveform_sig_rx =42;
26628: waveform_sig_rx =43;
26629: waveform_sig_rx =-165;
26630: waveform_sig_rx =29;
26631: waveform_sig_rx =148;
26632: waveform_sig_rx =-129;
26633: waveform_sig_rx =-23;
26634: waveform_sig_rx =216;
26635: waveform_sig_rx =-36;
26636: waveform_sig_rx =-70;
26637: waveform_sig_rx =255;
26638: waveform_sig_rx =29;
26639: waveform_sig_rx =-36;
26640: waveform_sig_rx =191;
26641: waveform_sig_rx =163;
26642: waveform_sig_rx =-34;
26643: waveform_sig_rx =119;
26644: waveform_sig_rx =243;
26645: waveform_sig_rx =10;
26646: waveform_sig_rx =34;
26647: waveform_sig_rx =326;
26648: waveform_sig_rx =70;
26649: waveform_sig_rx =59;
26650: waveform_sig_rx =238;
26651: waveform_sig_rx =93;
26652: waveform_sig_rx =212;
26653: waveform_sig_rx =146;
26654: waveform_sig_rx =248;
26655: waveform_sig_rx =-11;
26656: waveform_sig_rx =443;
26657: waveform_sig_rx =37;
26658: waveform_sig_rx =146;
26659: waveform_sig_rx =444;
26660: waveform_sig_rx =2;
26661: waveform_sig_rx =253;
26662: waveform_sig_rx =394;
26663: waveform_sig_rx =117;
26664: waveform_sig_rx =181;
26665: waveform_sig_rx =405;
26666: waveform_sig_rx =216;
26667: waveform_sig_rx =160;
26668: waveform_sig_rx =402;
26669: waveform_sig_rx =365;
26670: waveform_sig_rx =61;
26671: waveform_sig_rx =419;
26672: waveform_sig_rx =385;
26673: waveform_sig_rx =158;
26674: waveform_sig_rx =311;
26675: waveform_sig_rx =462;
26676: waveform_sig_rx =279;
26677: waveform_sig_rx =230;
26678: waveform_sig_rx =531;
26679: waveform_sig_rx =312;
26680: waveform_sig_rx =244;
26681: waveform_sig_rx =465;
26682: waveform_sig_rx =416;
26683: waveform_sig_rx =264;
26684: waveform_sig_rx =382;
26685: waveform_sig_rx =550;
26686: waveform_sig_rx =295;
26687: waveform_sig_rx =295;
26688: waveform_sig_rx =649;
26689: waveform_sig_rx =305;
26690: waveform_sig_rx =388;
26691: waveform_sig_rx =538;
26692: waveform_sig_rx =313;
26693: waveform_sig_rx =568;
26694: waveform_sig_rx =417;
26695: waveform_sig_rx =479;
26696: waveform_sig_rx =347;
26697: waveform_sig_rx =661;
26698: waveform_sig_rx =334;
26699: waveform_sig_rx =472;
26700: waveform_sig_rx =629;
26701: waveform_sig_rx =363;
26702: waveform_sig_rx =468;
26703: waveform_sig_rx =682;
26704: waveform_sig_rx =412;
26705: waveform_sig_rx =398;
26706: waveform_sig_rx =769;
26707: waveform_sig_rx =441;
26708: waveform_sig_rx =436;
26709: waveform_sig_rx =713;
26710: waveform_sig_rx =573;
26711: waveform_sig_rx =346;
26712: waveform_sig_rx =717;
26713: waveform_sig_rx =638;
26714: waveform_sig_rx =448;
26715: waveform_sig_rx =602;
26716: waveform_sig_rx =736;
26717: waveform_sig_rx =519;
26718: waveform_sig_rx =533;
26719: waveform_sig_rx =756;
26720: waveform_sig_rx =590;
26721: waveform_sig_rx =518;
26722: waveform_sig_rx =708;
26723: waveform_sig_rx =772;
26724: waveform_sig_rx =457;
26725: waveform_sig_rx =675;
26726: waveform_sig_rx =864;
26727: waveform_sig_rx =475;
26728: waveform_sig_rx =658;
26729: waveform_sig_rx =877;
26730: waveform_sig_rx =513;
26731: waveform_sig_rx =757;
26732: waveform_sig_rx =699;
26733: waveform_sig_rx =624;
26734: waveform_sig_rx =831;
26735: waveform_sig_rx =618;
26736: waveform_sig_rx =802;
26737: waveform_sig_rx =581;
26738: waveform_sig_rx =877;
26739: waveform_sig_rx =630;
26740: waveform_sig_rx =656;
26741: waveform_sig_rx =917;
26742: waveform_sig_rx =607;
26743: waveform_sig_rx =672;
26744: waveform_sig_rx =982;
26745: waveform_sig_rx =619;
26746: waveform_sig_rx =650;
26747: waveform_sig_rx =1014;
26748: waveform_sig_rx =646;
26749: waveform_sig_rx =688;
26750: waveform_sig_rx =968;
26751: waveform_sig_rx =780;
26752: waveform_sig_rx =603;
26753: waveform_sig_rx =965;
26754: waveform_sig_rx =814;
26755: waveform_sig_rx =711;
26756: waveform_sig_rx =826;
26757: waveform_sig_rx =917;
26758: waveform_sig_rx =774;
26759: waveform_sig_rx =725;
26760: waveform_sig_rx =988;
26761: waveform_sig_rx =859;
26762: waveform_sig_rx =690;
26763: waveform_sig_rx =985;
26764: waveform_sig_rx =957;
26765: waveform_sig_rx =626;
26766: waveform_sig_rx =1001;
26767: waveform_sig_rx =971;
26768: waveform_sig_rx =692;
26769: waveform_sig_rx =917;
26770: waveform_sig_rx =1012;
26771: waveform_sig_rx =810;
26772: waveform_sig_rx =899;
26773: waveform_sig_rx =881;
26774: waveform_sig_rx =907;
26775: waveform_sig_rx =949;
26776: waveform_sig_rx =863;
26777: waveform_sig_rx =997;
26778: waveform_sig_rx =746;
26779: waveform_sig_rx =1139;
26780: waveform_sig_rx =796;
26781: waveform_sig_rx =875;
26782: waveform_sig_rx =1139;
26783: waveform_sig_rx =789;
26784: waveform_sig_rx =904;
26785: waveform_sig_rx =1201;
26786: waveform_sig_rx =801;
26787: waveform_sig_rx =880;
26788: waveform_sig_rx =1273;
26789: waveform_sig_rx =772;
26790: waveform_sig_rx =948;
26791: waveform_sig_rx =1169;
26792: waveform_sig_rx =896;
26793: waveform_sig_rx =885;
26794: waveform_sig_rx =1108;
26795: waveform_sig_rx =1006;
26796: waveform_sig_rx =933;
26797: waveform_sig_rx =936;
26798: waveform_sig_rx =1168;
26799: waveform_sig_rx =905;
26800: waveform_sig_rx =885;
26801: waveform_sig_rx =1221;
26802: waveform_sig_rx =926;
26803: waveform_sig_rx =886;
26804: waveform_sig_rx =1180;
26805: waveform_sig_rx =1053;
26806: waveform_sig_rx =824;
26807: waveform_sig_rx =1136;
26808: waveform_sig_rx =1093;
26809: waveform_sig_rx =904;
26810: waveform_sig_rx =1046;
26811: waveform_sig_rx =1150;
26812: waveform_sig_rx =979;
26813: waveform_sig_rx =1029;
26814: waveform_sig_rx =1060;
26815: waveform_sig_rx =1087;
26816: waveform_sig_rx =1061;
26817: waveform_sig_rx =1059;
26818: waveform_sig_rx =1118;
26819: waveform_sig_rx =895;
26820: waveform_sig_rx =1327;
26821: waveform_sig_rx =883;
26822: waveform_sig_rx =1055;
26823: waveform_sig_rx =1291;
26824: waveform_sig_rx =848;
26825: waveform_sig_rx =1089;
26826: waveform_sig_rx =1310;
26827: waveform_sig_rx =881;
26828: waveform_sig_rx =1061;
26829: waveform_sig_rx =1342;
26830: waveform_sig_rx =881;
26831: waveform_sig_rx =1114;
26832: waveform_sig_rx =1223;
26833: waveform_sig_rx =1063;
26834: waveform_sig_rx =1016;
26835: waveform_sig_rx =1174;
26836: waveform_sig_rx =1177;
26837: waveform_sig_rx =999;
26838: waveform_sig_rx =1078;
26839: waveform_sig_rx =1330;
26840: waveform_sig_rx =953;
26841: waveform_sig_rx =1079;
26842: waveform_sig_rx =1329;
26843: waveform_sig_rx =1015;
26844: waveform_sig_rx =1048;
26845: waveform_sig_rx =1252;
26846: waveform_sig_rx =1145;
26847: waveform_sig_rx =984;
26848: waveform_sig_rx =1234;
26849: waveform_sig_rx =1222;
26850: waveform_sig_rx =1013;
26851: waveform_sig_rx =1124;
26852: waveform_sig_rx =1285;
26853: waveform_sig_rx =1043;
26854: waveform_sig_rx =1128;
26855: waveform_sig_rx =1182;
26856: waveform_sig_rx =1126;
26857: waveform_sig_rx =1154;
26858: waveform_sig_rx =1183;
26859: waveform_sig_rx =1129;
26860: waveform_sig_rx =1020;
26861: waveform_sig_rx =1406;
26862: waveform_sig_rx =916;
26863: waveform_sig_rx =1193;
26864: waveform_sig_rx =1313;
26865: waveform_sig_rx =926;
26866: waveform_sig_rx =1225;
26867: waveform_sig_rx =1298;
26868: waveform_sig_rx =962;
26869: waveform_sig_rx =1154;
26870: waveform_sig_rx =1342;
26871: waveform_sig_rx =985;
26872: waveform_sig_rx =1156;
26873: waveform_sig_rx =1279;
26874: waveform_sig_rx =1139;
26875: waveform_sig_rx =1009;
26876: waveform_sig_rx =1271;
26877: waveform_sig_rx =1221;
26878: waveform_sig_rx =1012;
26879: waveform_sig_rx =1160;
26880: waveform_sig_rx =1352;
26881: waveform_sig_rx =964;
26882: waveform_sig_rx =1172;
26883: waveform_sig_rx =1307;
26884: waveform_sig_rx =1038;
26885: waveform_sig_rx =1124;
26886: waveform_sig_rx =1224;
26887: waveform_sig_rx =1210;
26888: waveform_sig_rx =992;
26889: waveform_sig_rx =1205;
26890: waveform_sig_rx =1280;
26891: waveform_sig_rx =981;
26892: waveform_sig_rx =1170;
26893: waveform_sig_rx =1358;
26894: waveform_sig_rx =970;
26895: waveform_sig_rx =1199;
26896: waveform_sig_rx =1152;
26897: waveform_sig_rx =1101;
26898: waveform_sig_rx =1202;
26899: waveform_sig_rx =1154;
26900: waveform_sig_rx =1131;
26901: waveform_sig_rx =1071;
26902: waveform_sig_rx =1343;
26903: waveform_sig_rx =917;
26904: waveform_sig_rx =1204;
26905: waveform_sig_rx =1267;
26906: waveform_sig_rx =950;
26907: waveform_sig_rx =1221;
26908: waveform_sig_rx =1265;
26909: waveform_sig_rx =978;
26910: waveform_sig_rx =1132;
26911: waveform_sig_rx =1293;
26912: waveform_sig_rx =983;
26913: waveform_sig_rx =1095;
26914: waveform_sig_rx =1271;
26915: waveform_sig_rx =1118;
26916: waveform_sig_rx =933;
26917: waveform_sig_rx =1304;
26918: waveform_sig_rx =1121;
26919: waveform_sig_rx =973;
26920: waveform_sig_rx =1173;
26921: waveform_sig_rx =1241;
26922: waveform_sig_rx =972;
26923: waveform_sig_rx =1136;
26924: waveform_sig_rx =1238;
26925: waveform_sig_rx =1049;
26926: waveform_sig_rx =1018;
26927: waveform_sig_rx =1223;
26928: waveform_sig_rx =1169;
26929: waveform_sig_rx =903;
26930: waveform_sig_rx =1199;
26931: waveform_sig_rx =1198;
26932: waveform_sig_rx =898;
26933: waveform_sig_rx =1144;
26934: waveform_sig_rx =1244;
26935: waveform_sig_rx =902;
26936: waveform_sig_rx =1147;
26937: waveform_sig_rx =1041;
26938: waveform_sig_rx =1058;
26939: waveform_sig_rx =1117;
26940: waveform_sig_rx =1054;
26941: waveform_sig_rx =1039;
26942: waveform_sig_rx =983;
26943: waveform_sig_rx =1231;
26944: waveform_sig_rx =872;
26945: waveform_sig_rx =1112;
26946: waveform_sig_rx =1149;
26947: waveform_sig_rx =882;
26948: waveform_sig_rx =1079;
26949: waveform_sig_rx =1202;
26950: waveform_sig_rx =862;
26951: waveform_sig_rx =1006;
26952: waveform_sig_rx =1242;
26953: waveform_sig_rx =851;
26954: waveform_sig_rx =1000;
26955: waveform_sig_rx =1201;
26956: waveform_sig_rx =949;
26957: waveform_sig_rx =883;
26958: waveform_sig_rx =1213;
26959: waveform_sig_rx =941;
26960: waveform_sig_rx =932;
26961: waveform_sig_rx =1036;
26962: waveform_sig_rx =1117;
26963: waveform_sig_rx =867;
26964: waveform_sig_rx =955;
26965: waveform_sig_rx =1151;
26966: waveform_sig_rx =897;
26967: waveform_sig_rx =870;
26968: waveform_sig_rx =1131;
26969: waveform_sig_rx =1003;
26970: waveform_sig_rx =771;
26971: waveform_sig_rx =1135;
26972: waveform_sig_rx =1018;
26973: waveform_sig_rx =780;
26974: waveform_sig_rx =1032;
26975: waveform_sig_rx =1076;
26976: waveform_sig_rx =783;
26977: waveform_sig_rx =1052;
26978: waveform_sig_rx =881;
26979: waveform_sig_rx =978;
26980: waveform_sig_rx =962;
26981: waveform_sig_rx =894;
26982: waveform_sig_rx =946;
26983: waveform_sig_rx =831;
26984: waveform_sig_rx =1099;
26985: waveform_sig_rx =744;
26986: waveform_sig_rx =930;
26987: waveform_sig_rx =1060;
26988: waveform_sig_rx =692;
26989: waveform_sig_rx =916;
26990: waveform_sig_rx =1076;
26991: waveform_sig_rx =649;
26992: waveform_sig_rx =921;
26993: waveform_sig_rx =1076;
26994: waveform_sig_rx =637;
26995: waveform_sig_rx =906;
26996: waveform_sig_rx =983;
26997: waveform_sig_rx =765;
26998: waveform_sig_rx =729;
26999: waveform_sig_rx =994;
27000: waveform_sig_rx =798;
27001: waveform_sig_rx =757;
27002: waveform_sig_rx =844;
27003: waveform_sig_rx =941;
27004: waveform_sig_rx =683;
27005: waveform_sig_rx =768;
27006: waveform_sig_rx =963;
27007: waveform_sig_rx =700;
27008: waveform_sig_rx =679;
27009: waveform_sig_rx =988;
27010: waveform_sig_rx =735;
27011: waveform_sig_rx =596;
27012: waveform_sig_rx =943;
27013: waveform_sig_rx =770;
27014: waveform_sig_rx =637;
27015: waveform_sig_rx =810;
27016: waveform_sig_rx =854;
27017: waveform_sig_rx =617;
27018: waveform_sig_rx =799;
27019: waveform_sig_rx =676;
27020: waveform_sig_rx =776;
27021: waveform_sig_rx =695;
27022: waveform_sig_rx =754;
27023: waveform_sig_rx =715;
27024: waveform_sig_rx =610;
27025: waveform_sig_rx =937;
27026: waveform_sig_rx =477;
27027: waveform_sig_rx =757;
27028: waveform_sig_rx =838;
27029: waveform_sig_rx =431;
27030: waveform_sig_rx =784;
27031: waveform_sig_rx =832;
27032: waveform_sig_rx =409;
27033: waveform_sig_rx =746;
27034: waveform_sig_rx =836;
27035: waveform_sig_rx =431;
27036: waveform_sig_rx =715;
27037: waveform_sig_rx =740;
27038: waveform_sig_rx =543;
27039: waveform_sig_rx =520;
27040: waveform_sig_rx =737;
27041: waveform_sig_rx =588;
27042: waveform_sig_rx =508;
27043: waveform_sig_rx =566;
27044: waveform_sig_rx =758;
27045: waveform_sig_rx =392;
27046: waveform_sig_rx =568;
27047: waveform_sig_rx =767;
27048: waveform_sig_rx =384;
27049: waveform_sig_rx =527;
27050: waveform_sig_rx =720;
27051: waveform_sig_rx =475;
27052: waveform_sig_rx =451;
27053: waveform_sig_rx =627;
27054: waveform_sig_rx =567;
27055: waveform_sig_rx =386;
27056: waveform_sig_rx =518;
27057: waveform_sig_rx =667;
27058: waveform_sig_rx =328;
27059: waveform_sig_rx =585;
27060: waveform_sig_rx =449;
27061: waveform_sig_rx =508;
27062: waveform_sig_rx =455;
27063: waveform_sig_rx =508;
27064: waveform_sig_rx =418;
27065: waveform_sig_rx =383;
27066: waveform_sig_rx =671;
27067: waveform_sig_rx =194;
27068: waveform_sig_rx =535;
27069: waveform_sig_rx =549;
27070: waveform_sig_rx =144;
27071: waveform_sig_rx =577;
27072: waveform_sig_rx =488;
27073: waveform_sig_rx =141;
27074: waveform_sig_rx =535;
27075: waveform_sig_rx =469;
27076: waveform_sig_rx =222;
27077: waveform_sig_rx =424;
27078: waveform_sig_rx =439;
27079: waveform_sig_rx =330;
27080: waveform_sig_rx =184;
27081: waveform_sig_rx =505;
27082: waveform_sig_rx =307;
27083: waveform_sig_rx =195;
27084: waveform_sig_rx =375;
27085: waveform_sig_rx =428;
27086: waveform_sig_rx =112;
27087: waveform_sig_rx =343;
27088: waveform_sig_rx =426;
27089: waveform_sig_rx =127;
27090: waveform_sig_rx =252;
27091: waveform_sig_rx =382;
27092: waveform_sig_rx =205;
27093: waveform_sig_rx =142;
27094: waveform_sig_rx =345;
27095: waveform_sig_rx =305;
27096: waveform_sig_rx =83;
27097: waveform_sig_rx =259;
27098: waveform_sig_rx =389;
27099: waveform_sig_rx =15;
27100: waveform_sig_rx =308;
27101: waveform_sig_rx =128;
27102: waveform_sig_rx =203;
27103: waveform_sig_rx =175;
27104: waveform_sig_rx =238;
27105: waveform_sig_rx =82;
27106: waveform_sig_rx =142;
27107: waveform_sig_rx =329;
27108: waveform_sig_rx =-137;
27109: waveform_sig_rx =295;
27110: waveform_sig_rx =191;
27111: waveform_sig_rx =-108;
27112: waveform_sig_rx =279;
27113: waveform_sig_rx =144;
27114: waveform_sig_rx =-77;
27115: waveform_sig_rx =169;
27116: waveform_sig_rx =162;
27117: waveform_sig_rx =-31;
27118: waveform_sig_rx =50;
27119: waveform_sig_rx =221;
27120: waveform_sig_rx =-31;
27121: waveform_sig_rx =-126;
27122: waveform_sig_rx =281;
27123: waveform_sig_rx =-87;
27124: waveform_sig_rx =-61;
27125: waveform_sig_rx =90;
27126: waveform_sig_rx =94;
27127: waveform_sig_rx =-138;
27128: waveform_sig_rx =15;
27129: waveform_sig_rx =122;
27130: waveform_sig_rx =-171;
27131: waveform_sig_rx =-55;
27132: waveform_sig_rx =101;
27133: waveform_sig_rx =-94;
27134: waveform_sig_rx =-150;
27135: waveform_sig_rx =23;
27136: waveform_sig_rx =-2;
27137: waveform_sig_rx =-264;
27138: waveform_sig_rx =-25;
27139: waveform_sig_rx =74;
27140: waveform_sig_rx =-366;
27141: waveform_sig_rx =48;
27142: waveform_sig_rx =-215;
27143: waveform_sig_rx =-125;
27144: waveform_sig_rx =-98;
27145: waveform_sig_rx =-139;
27146: waveform_sig_rx =-204;
27147: waveform_sig_rx =-133;
27148: waveform_sig_rx =-34;
27149: waveform_sig_rx =-367;
27150: waveform_sig_rx =-58;
27151: waveform_sig_rx =-147;
27152: waveform_sig_rx =-364;
27153: waveform_sig_rx =-88;
27154: waveform_sig_rx =-100;
27155: waveform_sig_rx =-415;
27156: waveform_sig_rx =-139;
27157: waveform_sig_rx =-88;
27158: waveform_sig_rx =-402;
27159: waveform_sig_rx =-192;
27160: waveform_sig_rx =-105;
27161: waveform_sig_rx =-369;
27162: waveform_sig_rx =-370;
27163: waveform_sig_rx =-74;
27164: waveform_sig_rx =-377;
27165: waveform_sig_rx =-370;
27166: waveform_sig_rx =-234;
27167: waveform_sig_rx =-224;
27168: waveform_sig_rx =-472;
27169: waveform_sig_rx =-274;
27170: waveform_sig_rx =-223;
27171: waveform_sig_rx =-440;
27172: waveform_sig_rx =-384;
27173: waveform_sig_rx =-200;
27174: waveform_sig_rx =-379;
27175: waveform_sig_rx =-539;
27176: waveform_sig_rx =-183;
27177: waveform_sig_rx =-361;
27178: waveform_sig_rx =-586;
27179: waveform_sig_rx =-240;
27180: waveform_sig_rx =-330;
27181: waveform_sig_rx =-576;
27182: waveform_sig_rx =-259;
27183: waveform_sig_rx =-537;
27184: waveform_sig_rx =-320;
27185: waveform_sig_rx =-467;
27186: waveform_sig_rx =-415;
27187: waveform_sig_rx =-464;
27188: waveform_sig_rx =-479;
27189: waveform_sig_rx =-298;
27190: waveform_sig_rx =-674;
27191: waveform_sig_rx =-369;
27192: waveform_sig_rx =-364;
27193: waveform_sig_rx =-722;
27194: waveform_sig_rx =-351;
27195: waveform_sig_rx =-390;
27196: waveform_sig_rx =-740;
27197: waveform_sig_rx =-385;
27198: waveform_sig_rx =-399;
27199: waveform_sig_rx =-726;
27200: waveform_sig_rx =-471;
27201: waveform_sig_rx =-398;
27202: waveform_sig_rx =-682;
27203: waveform_sig_rx =-629;
27204: waveform_sig_rx =-356;
27205: waveform_sig_rx =-657;
27206: waveform_sig_rx =-612;
27207: waveform_sig_rx =-515;
27208: waveform_sig_rx =-506;
27209: waveform_sig_rx =-727;
27210: waveform_sig_rx =-591;
27211: waveform_sig_rx =-476;
27212: waveform_sig_rx =-756;
27213: waveform_sig_rx =-682;
27214: waveform_sig_rx =-408;
27215: waveform_sig_rx =-743;
27216: waveform_sig_rx =-763;
27217: waveform_sig_rx =-460;
27218: waveform_sig_rx =-730;
27219: waveform_sig_rx =-781;
27220: waveform_sig_rx =-569;
27221: waveform_sig_rx =-628;
27222: waveform_sig_rx =-793;
27223: waveform_sig_rx =-615;
27224: waveform_sig_rx =-769;
27225: waveform_sig_rx =-608;
27226: waveform_sig_rx =-786;
27227: waveform_sig_rx =-601;
27228: waveform_sig_rx =-800;
27229: waveform_sig_rx =-721;
27230: waveform_sig_rx =-563;
27231: waveform_sig_rx =-957;
27232: waveform_sig_rx =-586;
27233: waveform_sig_rx =-658;
27234: waveform_sig_rx =-961;
27235: waveform_sig_rx =-591;
27236: waveform_sig_rx =-664;
27237: waveform_sig_rx =-1005;
27238: waveform_sig_rx =-625;
27239: waveform_sig_rx =-649;
27240: waveform_sig_rx =-1006;
27241: waveform_sig_rx =-672;
27242: waveform_sig_rx =-693;
27243: waveform_sig_rx =-957;
27244: waveform_sig_rx =-810;
27245: waveform_sig_rx =-694;
27246: waveform_sig_rx =-871;
27247: waveform_sig_rx =-880;
27248: waveform_sig_rx =-801;
27249: waveform_sig_rx =-672;
27250: waveform_sig_rx =-1061;
27251: waveform_sig_rx =-755;
27252: waveform_sig_rx =-704;
27253: waveform_sig_rx =-1054;
27254: waveform_sig_rx =-837;
27255: waveform_sig_rx =-696;
27256: waveform_sig_rx =-962;
27257: waveform_sig_rx =-941;
27258: waveform_sig_rx =-712;
27259: waveform_sig_rx =-900;
27260: waveform_sig_rx =-1010;
27261: waveform_sig_rx =-783;
27262: waveform_sig_rx =-815;
27263: waveform_sig_rx =-1040;
27264: waveform_sig_rx =-825;
27265: waveform_sig_rx =-979;
27266: waveform_sig_rx =-824;
27267: waveform_sig_rx =-995;
27268: waveform_sig_rx =-805;
27269: waveform_sig_rx =-1057;
27270: waveform_sig_rx =-899;
27271: waveform_sig_rx =-805;
27272: waveform_sig_rx =-1199;
27273: waveform_sig_rx =-757;
27274: waveform_sig_rx =-904;
27275: waveform_sig_rx =-1188;
27276: waveform_sig_rx =-742;
27277: waveform_sig_rx =-943;
27278: waveform_sig_rx =-1206;
27279: waveform_sig_rx =-778;
27280: waveform_sig_rx =-946;
27281: waveform_sig_rx =-1171;
27282: waveform_sig_rx =-885;
27283: waveform_sig_rx =-931;
27284: waveform_sig_rx =-1087;
27285: waveform_sig_rx =-1069;
27286: waveform_sig_rx =-866;
27287: waveform_sig_rx =-1039;
27288: waveform_sig_rx =-1137;
27289: waveform_sig_rx =-912;
27290: waveform_sig_rx =-907;
27291: waveform_sig_rx =-1252;
27292: waveform_sig_rx =-875;
27293: waveform_sig_rx =-972;
27294: waveform_sig_rx =-1185;
27295: waveform_sig_rx =-984;
27296: waveform_sig_rx =-919;
27297: waveform_sig_rx =-1114;
27298: waveform_sig_rx =-1138;
27299: waveform_sig_rx =-888;
27300: waveform_sig_rx =-1046;
27301: waveform_sig_rx =-1199;
27302: waveform_sig_rx =-935;
27303: waveform_sig_rx =-977;
27304: waveform_sig_rx =-1222;
27305: waveform_sig_rx =-965;
27306: waveform_sig_rx =-1133;
27307: waveform_sig_rx =-1023;
27308: waveform_sig_rx =-1121;
27309: waveform_sig_rx =-974;
27310: waveform_sig_rx =-1247;
27311: waveform_sig_rx =-976;
27312: waveform_sig_rx =-1020;
27313: waveform_sig_rx =-1334;
27314: waveform_sig_rx =-895;
27315: waveform_sig_rx =-1142;
27316: waveform_sig_rx =-1278;
27317: waveform_sig_rx =-913;
27318: waveform_sig_rx =-1107;
27319: waveform_sig_rx =-1290;
27320: waveform_sig_rx =-971;
27321: waveform_sig_rx =-1090;
27322: waveform_sig_rx =-1278;
27323: waveform_sig_rx =-1039;
27324: waveform_sig_rx =-1035;
27325: waveform_sig_rx =-1229;
27326: waveform_sig_rx =-1189;
27327: waveform_sig_rx =-950;
27328: waveform_sig_rx =-1191;
27329: waveform_sig_rx =-1254;
27330: waveform_sig_rx =-983;
27331: waveform_sig_rx =-1099;
27332: waveform_sig_rx =-1336;
27333: waveform_sig_rx =-980;
27334: waveform_sig_rx =-1132;
27335: waveform_sig_rx =-1234;
27336: waveform_sig_rx =-1122;
27337: waveform_sig_rx =-1014;
27338: waveform_sig_rx =-1176;
27339: waveform_sig_rx =-1272;
27340: waveform_sig_rx =-941;
27341: waveform_sig_rx =-1171;
27342: waveform_sig_rx =-1311;
27343: waveform_sig_rx =-981;
27344: waveform_sig_rx =-1116;
27345: waveform_sig_rx =-1306;
27346: waveform_sig_rx =-1041;
27347: waveform_sig_rx =-1261;
27348: waveform_sig_rx =-1088;
27349: waveform_sig_rx =-1190;
27350: waveform_sig_rx =-1100;
27351: waveform_sig_rx =-1304;
27352: waveform_sig_rx =-1043;
27353: waveform_sig_rx =-1140;
27354: waveform_sig_rx =-1339;
27355: waveform_sig_rx =-975;
27356: waveform_sig_rx =-1203;
27357: waveform_sig_rx =-1284;
27358: waveform_sig_rx =-1019;
27359: waveform_sig_rx =-1126;
27360: waveform_sig_rx =-1370;
27361: waveform_sig_rx =-1029;
27362: waveform_sig_rx =-1104;
27363: waveform_sig_rx =-1338;
27364: waveform_sig_rx =-1063;
27365: waveform_sig_rx =-1047;
27366: waveform_sig_rx =-1310;
27367: waveform_sig_rx =-1186;
27368: waveform_sig_rx =-970;
27369: waveform_sig_rx =-1274;
27370: waveform_sig_rx =-1234;
27371: waveform_sig_rx =-1041;
27372: waveform_sig_rx =-1156;
27373: waveform_sig_rx =-1292;
27374: waveform_sig_rx =-1035;
27375: waveform_sig_rx =-1114;
27376: waveform_sig_rx =-1240;
27377: waveform_sig_rx =-1205;
27378: waveform_sig_rx =-978;
27379: waveform_sig_rx =-1242;
27380: waveform_sig_rx =-1275;
27381: waveform_sig_rx =-928;
27382: waveform_sig_rx =-1243;
27383: waveform_sig_rx =-1250;
27384: waveform_sig_rx =-989;
27385: waveform_sig_rx =-1151;
27386: waveform_sig_rx =-1265;
27387: waveform_sig_rx =-1057;
27388: waveform_sig_rx =-1254;
27389: waveform_sig_rx =-1069;
27390: waveform_sig_rx =-1201;
27391: waveform_sig_rx =-1077;
27392: waveform_sig_rx =-1272;
27393: waveform_sig_rx =-1033;
27394: waveform_sig_rx =-1137;
27395: waveform_sig_rx =-1273;
27396: waveform_sig_rx =-972;
27397: waveform_sig_rx =-1171;
27398: waveform_sig_rx =-1240;
27399: waveform_sig_rx =-1009;
27400: waveform_sig_rx =-1058;
27401: waveform_sig_rx =-1363;
27402: waveform_sig_rx =-945;
27403: waveform_sig_rx =-1038;
27404: waveform_sig_rx =-1362;
27405: waveform_sig_rx =-957;
27406: waveform_sig_rx =-1062;
27407: waveform_sig_rx =-1291;
27408: waveform_sig_rx =-1081;
27409: waveform_sig_rx =-1019;
27410: waveform_sig_rx =-1203;
27411: waveform_sig_rx =-1163;
27412: waveform_sig_rx =-1016;
27413: waveform_sig_rx =-1056;
27414: waveform_sig_rx =-1266;
27415: waveform_sig_rx =-989;
27416: waveform_sig_rx =-1029;
27417: waveform_sig_rx =-1230;
27418: waveform_sig_rx =-1089;
27419: waveform_sig_rx =-915;
27420: waveform_sig_rx =-1222;
27421: waveform_sig_rx =-1161;
27422: waveform_sig_rx =-872;
27423: waveform_sig_rx =-1204;
27424: waveform_sig_rx =-1168;
27425: waveform_sig_rx =-901;
27426: waveform_sig_rx =-1094;
27427: waveform_sig_rx =-1135;
27428: waveform_sig_rx =-983;
27429: waveform_sig_rx =-1168;
27430: waveform_sig_rx =-936;
27431: waveform_sig_rx =-1152;
27432: waveform_sig_rx =-940;
27433: waveform_sig_rx =-1169;
27434: waveform_sig_rx =-954;
27435: waveform_sig_rx =-975;
27436: waveform_sig_rx =-1223;
27437: waveform_sig_rx =-865;
27438: waveform_sig_rx =-1025;
27439: waveform_sig_rx =-1227;
27440: waveform_sig_rx =-810;
27441: waveform_sig_rx =-999;
27442: waveform_sig_rx =-1253;
27443: waveform_sig_rx =-765;
27444: waveform_sig_rx =-1019;
27445: waveform_sig_rx =-1183;
27446: waveform_sig_rx =-824;
27447: waveform_sig_rx =-956;
27448: waveform_sig_rx =-1130;
27449: waveform_sig_rx =-958;
27450: waveform_sig_rx =-863;
27451: waveform_sig_rx =-1039;
27452: waveform_sig_rx =-1042;
27453: waveform_sig_rx =-874;
27454: waveform_sig_rx =-935;
27455: waveform_sig_rx =-1153;
27456: waveform_sig_rx =-828;
27457: waveform_sig_rx =-894;
27458: waveform_sig_rx =-1108;
27459: waveform_sig_rx =-907;
27460: waveform_sig_rx =-774;
27461: waveform_sig_rx =-1084;
27462: waveform_sig_rx =-957;
27463: waveform_sig_rx =-730;
27464: waveform_sig_rx =-1042;
27465: waveform_sig_rx =-975;
27466: waveform_sig_rx =-808;
27467: waveform_sig_rx =-923;
27468: waveform_sig_rx =-986;
27469: waveform_sig_rx =-870;
27470: waveform_sig_rx =-956;
27471: waveform_sig_rx =-783;
27472: waveform_sig_rx =-1007;
27473: waveform_sig_rx =-739;
27474: waveform_sig_rx =-1063;
27475: waveform_sig_rx =-739;
27476: waveform_sig_rx =-824;
27477: waveform_sig_rx =-1088;
27478: waveform_sig_rx =-618;
27479: waveform_sig_rx =-923;
27480: waveform_sig_rx =-1027;
27481: waveform_sig_rx =-588;
27482: waveform_sig_rx =-927;
27483: waveform_sig_rx =-1005;
27484: waveform_sig_rx =-608;
27485: waveform_sig_rx =-867;
27486: waveform_sig_rx =-950;
27487: waveform_sig_rx =-694;
27488: waveform_sig_rx =-753;
27489: waveform_sig_rx =-946;
27490: waveform_sig_rx =-765;
27491: waveform_sig_rx =-667;
27492: waveform_sig_rx =-866;
27493: waveform_sig_rx =-846;
27494: waveform_sig_rx =-669;
27495: waveform_sig_rx =-741;
27496: waveform_sig_rx =-951;
27497: waveform_sig_rx =-596;
27498: waveform_sig_rx =-725;
27499: waveform_sig_rx =-933;
27500: waveform_sig_rx =-629;
27501: waveform_sig_rx =-656;
27502: waveform_sig_rx =-875;
27503: waveform_sig_rx =-715;
27504: waveform_sig_rx =-618;
27505: waveform_sig_rx =-765;
27506: waveform_sig_rx =-821;
27507: waveform_sig_rx =-576;
27508: waveform_sig_rx =-675;
27509: waveform_sig_rx =-828;
27510: waveform_sig_rx =-588;
27511: waveform_sig_rx =-769;
27512: waveform_sig_rx =-615;
27513: waveform_sig_rx =-714;
27514: waveform_sig_rx =-562;
27515: waveform_sig_rx =-852;
27516: waveform_sig_rx =-466;
27517: waveform_sig_rx =-680;
27518: waveform_sig_rx =-811;
27519: waveform_sig_rx =-401;
27520: waveform_sig_rx =-747;
27521: waveform_sig_rx =-750;
27522: waveform_sig_rx =-386;
27523: waveform_sig_rx =-713;
27524: waveform_sig_rx =-741;
27525: waveform_sig_rx =-377;
27526: waveform_sig_rx =-658;
27527: waveform_sig_rx =-653;
27528: waveform_sig_rx =-485;
27529: waveform_sig_rx =-492;
27530: waveform_sig_rx =-694;
27531: waveform_sig_rx =-557;
27532: waveform_sig_rx =-394;
27533: waveform_sig_rx =-653;
27534: waveform_sig_rx =-600;
27535: waveform_sig_rx =-366;
27536: waveform_sig_rx =-557;
27537: waveform_sig_rx =-660;
27538: waveform_sig_rx =-331;
27539: waveform_sig_rx =-511;
27540: waveform_sig_rx =-621;
27541: waveform_sig_rx =-428;
27542: waveform_sig_rx =-391;
27543: waveform_sig_rx =-611;
27544: waveform_sig_rx =-513;
27545: waveform_sig_rx =-314;
27546: waveform_sig_rx =-525;
27547: waveform_sig_rx =-595;
27548: waveform_sig_rx =-265;
27549: waveform_sig_rx =-473;
27550: waveform_sig_rx =-559;
27551: waveform_sig_rx =-283;
27552: waveform_sig_rx =-541;
27553: waveform_sig_rx =-321;
27554: waveform_sig_rx =-445;
27555: waveform_sig_rx =-327;
27556: waveform_sig_rx =-564;
27557: waveform_sig_rx =-208;
27558: waveform_sig_rx =-443;
27559: waveform_sig_rx =-515;
27560: waveform_sig_rx =-141;
27561: waveform_sig_rx =-484;
27562: waveform_sig_rx =-448;
27563: waveform_sig_rx =-123;
27564: waveform_sig_rx =-438;
27565: waveform_sig_rx =-450;
27566: waveform_sig_rx =-147;
27567: waveform_sig_rx =-361;
27568: waveform_sig_rx =-410;
27569: waveform_sig_rx =-233;
27570: waveform_sig_rx =-196;
27571: waveform_sig_rx =-509;
27572: waveform_sig_rx =-235;
27573: waveform_sig_rx =-123;
27574: waveform_sig_rx =-457;
27575: waveform_sig_rx =-265;
27576: waveform_sig_rx =-133;
27577: waveform_sig_rx =-293;
27578: waveform_sig_rx =-339;
27579: waveform_sig_rx =-108;
27580: waveform_sig_rx =-208;
27581: waveform_sig_rx =-354;
27582: waveform_sig_rx =-152;
27583: waveform_sig_rx =-79;
27584: waveform_sig_rx =-340;
27585: waveform_sig_rx =-229;
27586: waveform_sig_rx =-20;
27587: waveform_sig_rx =-263;
27588: waveform_sig_rx =-277;
27589: waveform_sig_rx =46;
27590: waveform_sig_rx =-224;
27591: waveform_sig_rx =-240;
27592: waveform_sig_rx =-15;
27593: waveform_sig_rx =-287;
27594: waveform_sig_rx =-10;
27595: waveform_sig_rx =-179;
27596: waveform_sig_rx =-56;
27597: waveform_sig_rx =-231;
27598: waveform_sig_rx =69;
27599: waveform_sig_rx =-154;
27600: waveform_sig_rx =-164;
27601: waveform_sig_rx =113;
27602: waveform_sig_rx =-162;
27603: waveform_sig_rx =-164;
27604: waveform_sig_rx =131;
27605: waveform_sig_rx =-113;
27606: waveform_sig_rx =-221;
27607: waveform_sig_rx =189;
27608: waveform_sig_rx =-82;
27609: waveform_sig_rx =-157;
27610: waveform_sig_rx =115;
27611: waveform_sig_rx =64;
27612: waveform_sig_rx =-209;
27613: waveform_sig_rx =101;
27614: waveform_sig_rx =121;
27615: waveform_sig_rx =-114;
27616: waveform_sig_rx =33;
27617: waveform_sig_rx =151;
27618: waveform_sig_rx =23;
27619: waveform_sig_rx =-56;
27620: waveform_sig_rx =203;
27621: waveform_sig_rx =85;
27622: waveform_sig_rx =-76;
27623: waveform_sig_rx =161;
27624: waveform_sig_rx =233;
27625: waveform_sig_rx =-72;
27626: waveform_sig_rx =92;
27627: waveform_sig_rx =299;
27628: waveform_sig_rx =-35;
27629: waveform_sig_rx =62;
27630: waveform_sig_rx =347;
27631: waveform_sig_rx =8;
27632: waveform_sig_rx =151;
27633: waveform_sig_rx =201;
27634: waveform_sig_rx =50;
27635: waveform_sig_rx =314;
27636: waveform_sig_rx =49;
27637: waveform_sig_rx =309;
27638: waveform_sig_rx =30;
27639: waveform_sig_rx =326;
27640: waveform_sig_rx =191;
27641: waveform_sig_rx =59;
27642: waveform_sig_rx =428;
27643: waveform_sig_rx =127;
27644: waveform_sig_rx =105;
27645: waveform_sig_rx =513;
27646: waveform_sig_rx =124;
27647: waveform_sig_rx =123;
27648: waveform_sig_rx =489;
27649: waveform_sig_rx =176;
27650: waveform_sig_rx =164;
27651: waveform_sig_rx =407;
27652: waveform_sig_rx =340;
27653: waveform_sig_rx =84;
27654: waveform_sig_rx =438;
27655: waveform_sig_rx =364;
27656: waveform_sig_rx =209;
27657: waveform_sig_rx =347;
27658: waveform_sig_rx =399;
27659: waveform_sig_rx =335;
27660: waveform_sig_rx =187;
27661: waveform_sig_rx =490;
27662: waveform_sig_rx =385;
27663: waveform_sig_rx =143;
27664: waveform_sig_rx =491;
27665: waveform_sig_rx =464;
27666: waveform_sig_rx =163;
27667: waveform_sig_rx =454;
27668: waveform_sig_rx =507;
27669: waveform_sig_rx =276;
27670: waveform_sig_rx =379;
27671: waveform_sig_rx =556;
27672: waveform_sig_rx =368;
27673: waveform_sig_rx =397;
27674: waveform_sig_rx =452;
27675: waveform_sig_rx =396;
27676: waveform_sig_rx =543;
27677: waveform_sig_rx =373;
27678: waveform_sig_rx =595;
27679: waveform_sig_rx =250;
27680: waveform_sig_rx =672;
27681: waveform_sig_rx =413;
27682: waveform_sig_rx =339;
27683: waveform_sig_rx =755;
27684: waveform_sig_rx =351;
27685: waveform_sig_rx =420;
27686: waveform_sig_rx =785;
27687: waveform_sig_rx =365;
27688: waveform_sig_rx =408;
27689: waveform_sig_rx =760;
27690: waveform_sig_rx =410;
27691: waveform_sig_rx =450;
27692: waveform_sig_rx =691;
27693: waveform_sig_rx =545;
27694: waveform_sig_rx =388;
27695: waveform_sig_rx =667;
27696: waveform_sig_rx =625;
27697: waveform_sig_rx =511;
27698: waveform_sig_rx =524;
27699: waveform_sig_rx =719;
27700: waveform_sig_rx =589;
27701: waveform_sig_rx =418;
27702: waveform_sig_rx =850;
27703: waveform_sig_rx =574;
27704: waveform_sig_rx =451;
27705: waveform_sig_rx =781;
27706: waveform_sig_rx =665;
27707: waveform_sig_rx =521;
27708: waveform_sig_rx =695;
27709: waveform_sig_rx =756;
27710: waveform_sig_rx =560;
27711: waveform_sig_rx =592;
27712: waveform_sig_rx =857;
27713: waveform_sig_rx =608;
27714: waveform_sig_rx =623;
27715: waveform_sig_rx =749;
27716: waveform_sig_rx =634;
27717: waveform_sig_rx =767;
27718: waveform_sig_rx =645;
27719: waveform_sig_rx =797;
27720: waveform_sig_rx =508;
27721: waveform_sig_rx =943;
27722: waveform_sig_rx =611;
27723: waveform_sig_rx =603;
27724: waveform_sig_rx =974;
27725: waveform_sig_rx =549;
27726: waveform_sig_rx =685;
27727: waveform_sig_rx =1021;
27728: waveform_sig_rx =567;
27729: waveform_sig_rx =711;
27730: waveform_sig_rx =994;
27731: waveform_sig_rx =616;
27732: waveform_sig_rx =739;
27733: waveform_sig_rx =867;
27734: waveform_sig_rx =821;
27735: waveform_sig_rx =640;
27736: waveform_sig_rx =865;
27737: waveform_sig_rx =915;
27738: waveform_sig_rx =681;
27739: waveform_sig_rx =763;
27740: waveform_sig_rx =1007;
27741: waveform_sig_rx =721;
27742: waveform_sig_rx =730;
27743: waveform_sig_rx =1026;
27744: waveform_sig_rx =762;
27745: waveform_sig_rx =745;
27746: waveform_sig_rx =961;
27747: waveform_sig_rx =912;
27748: waveform_sig_rx =721;
27749: waveform_sig_rx =875;
27750: waveform_sig_rx =989;
27751: waveform_sig_rx =748;
27752: waveform_sig_rx =813;
27753: waveform_sig_rx =1059;
27754: waveform_sig_rx =792;
27755: waveform_sig_rx =857;
27756: waveform_sig_rx =956;
27757: waveform_sig_rx =849;
27758: waveform_sig_rx =940;
27759: waveform_sig_rx =899;
27760: waveform_sig_rx =945;
27761: waveform_sig_rx =742;
27762: waveform_sig_rx =1168;
27763: waveform_sig_rx =741;
27764: waveform_sig_rx =904;
27765: waveform_sig_rx =1152;
27766: waveform_sig_rx =724;
27767: waveform_sig_rx =962;
27768: waveform_sig_rx =1134;
27769: waveform_sig_rx =801;
27770: waveform_sig_rx =904;
27771: waveform_sig_rx =1164;
27772: waveform_sig_rx =866;
27773: waveform_sig_rx =913;
27774: waveform_sig_rx =1076;
27775: waveform_sig_rx =1014;
27776: waveform_sig_rx =799;
27777: waveform_sig_rx =1102;
27778: waveform_sig_rx =1091;
27779: waveform_sig_rx =839;
27780: waveform_sig_rx =1004;
27781: waveform_sig_rx =1162;
27782: waveform_sig_rx =870;
27783: waveform_sig_rx =978;
27784: waveform_sig_rx =1161;
27785: waveform_sig_rx =950;
27786: waveform_sig_rx =931;
27787: waveform_sig_rx =1098;
27788: waveform_sig_rx =1097;
27789: waveform_sig_rx =861;
27790: waveform_sig_rx =1065;
27791: waveform_sig_rx =1191;
27792: waveform_sig_rx =867;
27793: waveform_sig_rx =1003;
27794: waveform_sig_rx =1253;
27795: waveform_sig_rx =904;
27796: waveform_sig_rx =1055;
27797: waveform_sig_rx =1074;
27798: waveform_sig_rx =982;
27799: waveform_sig_rx =1119;
27800: waveform_sig_rx =1049;
27801: waveform_sig_rx =1081;
27802: waveform_sig_rx =926;
27803: waveform_sig_rx =1282;
27804: waveform_sig_rx =874;
27805: waveform_sig_rx =1079;
27806: waveform_sig_rx =1218;
27807: waveform_sig_rx =908;
27808: waveform_sig_rx =1086;
27809: waveform_sig_rx =1215;
27810: waveform_sig_rx =962;
27811: waveform_sig_rx =979;
27812: waveform_sig_rx =1287;
27813: waveform_sig_rx =981;
27814: waveform_sig_rx =1000;
27815: waveform_sig_rx =1270;
27816: waveform_sig_rx =1094;
27817: waveform_sig_rx =900;
27818: waveform_sig_rx =1254;
27819: waveform_sig_rx =1129;
27820: waveform_sig_rx =975;
27821: waveform_sig_rx =1126;
27822: waveform_sig_rx =1247;
27823: waveform_sig_rx =995;
27824: waveform_sig_rx =1079;
27825: waveform_sig_rx =1261;
27826: waveform_sig_rx =1079;
27827: waveform_sig_rx =1012;
27828: waveform_sig_rx =1217;
27829: waveform_sig_rx =1239;
27830: waveform_sig_rx =915;
27831: waveform_sig_rx =1200;
27832: waveform_sig_rx =1254;
27833: waveform_sig_rx =921;
27834: waveform_sig_rx =1150;
27835: waveform_sig_rx =1294;
27836: waveform_sig_rx =968;
27837: waveform_sig_rx =1200;
27838: waveform_sig_rx =1107;
27839: waveform_sig_rx =1120;
27840: waveform_sig_rx =1201;
27841: waveform_sig_rx =1104;
27842: waveform_sig_rx =1188;
27843: waveform_sig_rx =992;
27844: waveform_sig_rx =1330;
27845: waveform_sig_rx =961;
27846: waveform_sig_rx =1129;
27847: waveform_sig_rx =1266;
27848: waveform_sig_rx =965;
27849: waveform_sig_rx =1123;
27850: waveform_sig_rx =1307;
27851: waveform_sig_rx =1011;
27852: waveform_sig_rx =1030;
27853: waveform_sig_rx =1398;
27854: waveform_sig_rx =983;
27855: waveform_sig_rx =1056;
27856: waveform_sig_rx =1360;
27857: waveform_sig_rx =1048;
27858: waveform_sig_rx =1011;
27859: waveform_sig_rx =1311;
27860: waveform_sig_rx =1128;
27861: waveform_sig_rx =1105;
27862: waveform_sig_rx =1116;
27863: waveform_sig_rx =1295;
27864: waveform_sig_rx =1042;
27865: waveform_sig_rx =1076;
27866: waveform_sig_rx =1339;
27867: waveform_sig_rx =1075;
27868: waveform_sig_rx =1064;
27869: waveform_sig_rx =1285;
27870: waveform_sig_rx =1212;
27871: waveform_sig_rx =951;
27872: waveform_sig_rx =1242;
27873: waveform_sig_rx =1269;
27874: waveform_sig_rx =958;
27875: waveform_sig_rx =1199;
27876: waveform_sig_rx =1277;
27877: waveform_sig_rx =1008;
27878: waveform_sig_rx =1211;
27879: waveform_sig_rx =1082;
27880: waveform_sig_rx =1173;
27881: waveform_sig_rx =1159;
27882: waveform_sig_rx =1087;
27883: waveform_sig_rx =1208;
27884: waveform_sig_rx =974;
27885: waveform_sig_rx =1363;
27886: waveform_sig_rx =983;
27887: waveform_sig_rx =1096;
27888: waveform_sig_rx =1334;
27889: waveform_sig_rx =932;
27890: waveform_sig_rx =1117;
27891: waveform_sig_rx =1362;
27892: waveform_sig_rx =904;
27893: waveform_sig_rx =1081;
27894: waveform_sig_rx =1372;
27895: waveform_sig_rx =898;
27896: waveform_sig_rx =1131;
27897: waveform_sig_rx =1258;
27898: waveform_sig_rx =1059;
27899: waveform_sig_rx =1012;
27900: waveform_sig_rx =1228;
27901: waveform_sig_rx =1146;
27902: waveform_sig_rx =1015;
27903: waveform_sig_rx =1094;
27904: waveform_sig_rx =1297;
27905: waveform_sig_rx =948;
27906: waveform_sig_rx =1063;
27907: waveform_sig_rx =1266;
27908: waveform_sig_rx =1018;
27909: waveform_sig_rx =1005;
27910: waveform_sig_rx =1252;
27911: waveform_sig_rx =1137;
27912: waveform_sig_rx =903;
27913: waveform_sig_rx =1228;
27914: waveform_sig_rx =1146;
27915: waveform_sig_rx =950;
27916: waveform_sig_rx =1138;
27917: waveform_sig_rx =1176;
27918: waveform_sig_rx =995;
27919: waveform_sig_rx =1075;
27920: waveform_sig_rx =1054;
27921: waveform_sig_rx =1125;
27922: waveform_sig_rx =1033;
27923: waveform_sig_rx =1098;
27924: waveform_sig_rx =1093;
27925: waveform_sig_rx =899;
27926: waveform_sig_rx =1334;
27927: waveform_sig_rx =835;
27928: waveform_sig_rx =1065;
27929: waveform_sig_rx =1244;
27930: waveform_sig_rx =771;
27931: waveform_sig_rx =1106;
27932: waveform_sig_rx =1199;
27933: waveform_sig_rx =815;
27934: waveform_sig_rx =1047;
27935: waveform_sig_rx =1198;
27936: waveform_sig_rx =849;
27937: waveform_sig_rx =1036;
27938: waveform_sig_rx =1128;
27939: waveform_sig_rx =984;
27940: waveform_sig_rx =881;
27941: waveform_sig_rx =1162;
27942: waveform_sig_rx =1023;
27943: waveform_sig_rx =895;
27944: waveform_sig_rx =998;
27945: waveform_sig_rx =1167;
27946: waveform_sig_rx =850;
27947: waveform_sig_rx =965;
27948: waveform_sig_rx =1168;
27949: waveform_sig_rx =861;
27950: waveform_sig_rx =915;
27951: waveform_sig_rx =1141;
27952: waveform_sig_rx =945;
27953: waveform_sig_rx =860;
27954: waveform_sig_rx =1070;
27955: waveform_sig_rx =1012;
27956: waveform_sig_rx =874;
27957: waveform_sig_rx =952;
27958: waveform_sig_rx =1131;
27959: waveform_sig_rx =833;
27960: waveform_sig_rx =934;
27961: waveform_sig_rx =975;
27962: waveform_sig_rx =916;
27963: waveform_sig_rx =934;
27964: waveform_sig_rx =983;
27965: waveform_sig_rx =858;
27966: waveform_sig_rx =855;
27967: waveform_sig_rx =1143;
27968: waveform_sig_rx =658;
27969: waveform_sig_rx =1012;
27970: waveform_sig_rx =1006;
27971: waveform_sig_rx =677;
27972: waveform_sig_rx =961;
27973: waveform_sig_rx =1028;
27974: waveform_sig_rx =666;
27975: waveform_sig_rx =891;
27976: waveform_sig_rx =1047;
27977: waveform_sig_rx =672;
27978: waveform_sig_rx =899;
27979: waveform_sig_rx =959;
27980: waveform_sig_rx =823;
27981: waveform_sig_rx =722;
27982: waveform_sig_rx =984;
27983: waveform_sig_rx =875;
27984: waveform_sig_rx =683;
27985: waveform_sig_rx =855;
27986: waveform_sig_rx =993;
27987: waveform_sig_rx =608;
27988: waveform_sig_rx =870;
27989: waveform_sig_rx =936;
27990: waveform_sig_rx =687;
27991: waveform_sig_rx =783;
27992: waveform_sig_rx =865;
27993: waveform_sig_rx =832;
27994: waveform_sig_rx =640;
27995: waveform_sig_rx =856;
27996: waveform_sig_rx =902;
27997: waveform_sig_rx =579;
27998: waveform_sig_rx =807;
27999: waveform_sig_rx =949;
28000: waveform_sig_rx =557;
28001: waveform_sig_rx =835;
28002: waveform_sig_rx =705;
28003: waveform_sig_rx =718;
28004: waveform_sig_rx =760;
28005: waveform_sig_rx =725;
28006: waveform_sig_rx =685;
28007: waveform_sig_rx =643;
28008: waveform_sig_rx =874;
28009: waveform_sig_rx =469;
28010: waveform_sig_rx =755;
28011: waveform_sig_rx =783;
28012: waveform_sig_rx =471;
28013: waveform_sig_rx =762;
28014: waveform_sig_rx =787;
28015: waveform_sig_rx =473;
28016: waveform_sig_rx =710;
28017: waveform_sig_rx =795;
28018: waveform_sig_rx =516;
28019: waveform_sig_rx =636;
28020: waveform_sig_rx =759;
28021: waveform_sig_rx =612;
28022: waveform_sig_rx =428;
28023: waveform_sig_rx =847;
28024: waveform_sig_rx =578;
28025: waveform_sig_rx =470;
28026: waveform_sig_rx =699;
28027: waveform_sig_rx =678;
28028: waveform_sig_rx =449;
28029: waveform_sig_rx =612;
28030: waveform_sig_rx =688;
28031: waveform_sig_rx =510;
28032: waveform_sig_rx =479;
28033: waveform_sig_rx =684;
28034: waveform_sig_rx =586;
28035: waveform_sig_rx =358;
28036: waveform_sig_rx =679;
28037: waveform_sig_rx =601;
28038: waveform_sig_rx =324;
28039: waveform_sig_rx =584;
28040: waveform_sig_rx =648;
28041: waveform_sig_rx =305;
28042: waveform_sig_rx =598;
28043: waveform_sig_rx =422;
28044: waveform_sig_rx =487;
28045: waveform_sig_rx =517;
28046: waveform_sig_rx =480;
28047: waveform_sig_rx =437;
28048: waveform_sig_rx =420;
28049: waveform_sig_rx =624;
28050: waveform_sig_rx =245;
28051: waveform_sig_rx =530;
28052: waveform_sig_rx =512;
28053: waveform_sig_rx =243;
28054: waveform_sig_rx =466;
28055: waveform_sig_rx =545;
28056: waveform_sig_rx =235;
28057: waveform_sig_rx =387;
28058: waveform_sig_rx =559;
28059: waveform_sig_rx =202;
28060: waveform_sig_rx =345;
28061: waveform_sig_rx =542;
28062: waveform_sig_rx =251;
28063: waveform_sig_rx =203;
28064: waveform_sig_rx =580;
28065: waveform_sig_rx =215;
28066: waveform_sig_rx =253;
28067: waveform_sig_rx =354;
28068: waveform_sig_rx =392;
28069: waveform_sig_rx =201;
28070: waveform_sig_rx =271;
28071: waveform_sig_rx =443;
28072: waveform_sig_rx =199;
28073: waveform_sig_rx =167;
28074: waveform_sig_rx =462;
28075: waveform_sig_rx =231;
28076: waveform_sig_rx =87;
28077: waveform_sig_rx =407;
28078: waveform_sig_rx =283;
28079: waveform_sig_rx =66;
28080: waveform_sig_rx =322;
28081: waveform_sig_rx =339;
28082: waveform_sig_rx =36;
28083: waveform_sig_rx =349;
28084: waveform_sig_rx =90;
28085: waveform_sig_rx =252;
28086: waveform_sig_rx =200;
28087: waveform_sig_rx =150;
28088: waveform_sig_rx =171;
28089: waveform_sig_rx =77;
28090: waveform_sig_rx =326;
28091: waveform_sig_rx =-51;
28092: waveform_sig_rx =175;
28093: waveform_sig_rx =274;
28094: waveform_sig_rx =-80;
28095: waveform_sig_rx =180;
28096: waveform_sig_rx =303;
28097: waveform_sig_rx =-148;
28098: waveform_sig_rx =179;
28099: waveform_sig_rx =260;
28100: waveform_sig_rx =-150;
28101: waveform_sig_rx =127;
28102: waveform_sig_rx =196;
28103: waveform_sig_rx =-47;
28104: waveform_sig_rx =-56;
28105: waveform_sig_rx =246;
28106: waveform_sig_rx =-43;
28107: waveform_sig_rx =-29;
28108: waveform_sig_rx =47;
28109: waveform_sig_rx =108;
28110: waveform_sig_rx =-98;
28111: waveform_sig_rx =-43;
28112: waveform_sig_rx =184;
28113: waveform_sig_rx =-134;
28114: waveform_sig_rx =-120;
28115: waveform_sig_rx =208;
28116: waveform_sig_rx =-131;
28117: waveform_sig_rx =-193;
28118: waveform_sig_rx =111;
28119: waveform_sig_rx =-108;
28120: waveform_sig_rx =-185;
28121: waveform_sig_rx =-14;
28122: waveform_sig_rx =7;
28123: waveform_sig_rx =-242;
28124: waveform_sig_rx =-30;
28125: waveform_sig_rx =-187;
28126: waveform_sig_rx =-43;
28127: waveform_sig_rx =-154;
28128: waveform_sig_rx =-97;
28129: waveform_sig_rx =-170;
28130: waveform_sig_rx =-244;
28131: waveform_sig_rx =53;
28132: waveform_sig_rx =-388;
28133: waveform_sig_rx =-104;
28134: waveform_sig_rx =-16;
28135: waveform_sig_rx =-450;
28136: waveform_sig_rx =-57;
28137: waveform_sig_rx =-51;
28138: waveform_sig_rx =-498;
28139: waveform_sig_rx =-75;
28140: waveform_sig_rx =-113;
28141: waveform_sig_rx =-439;
28142: waveform_sig_rx =-139;
28143: waveform_sig_rx =-167;
28144: waveform_sig_rx =-320;
28145: waveform_sig_rx =-374;
28146: waveform_sig_rx =-102;
28147: waveform_sig_rx =-324;
28148: waveform_sig_rx =-365;
28149: waveform_sig_rx =-259;
28150: waveform_sig_rx =-172;
28151: waveform_sig_rx =-469;
28152: waveform_sig_rx =-298;
28153: waveform_sig_rx =-138;
28154: waveform_sig_rx =-491;
28155: waveform_sig_rx =-366;
28156: waveform_sig_rx =-129;
28157: waveform_sig_rx =-459;
28158: waveform_sig_rx =-418;
28159: waveform_sig_rx =-233;
28160: waveform_sig_rx =-374;
28161: waveform_sig_rx =-469;
28162: waveform_sig_rx =-355;
28163: waveform_sig_rx =-236;
28164: waveform_sig_rx =-566;
28165: waveform_sig_rx =-347;
28166: waveform_sig_rx =-450;
28167: waveform_sig_rx =-377;
28168: waveform_sig_rx =-456;
28169: waveform_sig_rx =-369;
28170: waveform_sig_rx =-536;
28171: waveform_sig_rx =-474;
28172: waveform_sig_rx =-281;
28173: waveform_sig_rx =-734;
28174: waveform_sig_rx =-326;
28175: waveform_sig_rx =-380;
28176: waveform_sig_rx =-741;
28177: waveform_sig_rx =-295;
28178: waveform_sig_rx =-408;
28179: waveform_sig_rx =-752;
28180: waveform_sig_rx =-366;
28181: waveform_sig_rx =-452;
28182: waveform_sig_rx =-683;
28183: waveform_sig_rx =-466;
28184: waveform_sig_rx =-460;
28185: waveform_sig_rx =-577;
28186: waveform_sig_rx =-670;
28187: waveform_sig_rx =-364;
28188: waveform_sig_rx =-593;
28189: waveform_sig_rx =-704;
28190: waveform_sig_rx =-492;
28191: waveform_sig_rx =-458;
28192: waveform_sig_rx =-773;
28193: waveform_sig_rx =-512;
28194: waveform_sig_rx =-462;
28195: waveform_sig_rx =-771;
28196: waveform_sig_rx =-624;
28197: waveform_sig_rx =-479;
28198: waveform_sig_rx =-698;
28199: waveform_sig_rx =-722;
28200: waveform_sig_rx =-542;
28201: waveform_sig_rx =-613;
28202: waveform_sig_rx =-799;
28203: waveform_sig_rx =-614;
28204: waveform_sig_rx =-525;
28205: waveform_sig_rx =-859;
28206: waveform_sig_rx =-582;
28207: waveform_sig_rx =-715;
28208: waveform_sig_rx =-667;
28209: waveform_sig_rx =-720;
28210: waveform_sig_rx =-615;
28211: waveform_sig_rx =-834;
28212: waveform_sig_rx =-668;
28213: waveform_sig_rx =-587;
28214: waveform_sig_rx =-977;
28215: waveform_sig_rx =-512;
28216: waveform_sig_rx =-731;
28217: waveform_sig_rx =-930;
28218: waveform_sig_rx =-560;
28219: waveform_sig_rx =-735;
28220: waveform_sig_rx =-923;
28221: waveform_sig_rx =-683;
28222: waveform_sig_rx =-677;
28223: waveform_sig_rx =-916;
28224: waveform_sig_rx =-767;
28225: waveform_sig_rx =-663;
28226: waveform_sig_rx =-896;
28227: waveform_sig_rx =-932;
28228: waveform_sig_rx =-595;
28229: waveform_sig_rx =-885;
28230: waveform_sig_rx =-929;
28231: waveform_sig_rx =-716;
28232: waveform_sig_rx =-741;
28233: waveform_sig_rx =-1009;
28234: waveform_sig_rx =-730;
28235: waveform_sig_rx =-759;
28236: waveform_sig_rx =-978;
28237: waveform_sig_rx =-856;
28238: waveform_sig_rx =-746;
28239: waveform_sig_rx =-882;
28240: waveform_sig_rx =-1012;
28241: waveform_sig_rx =-722;
28242: waveform_sig_rx =-834;
28243: waveform_sig_rx =-1095;
28244: waveform_sig_rx =-757;
28245: waveform_sig_rx =-794;
28246: waveform_sig_rx =-1107;
28247: waveform_sig_rx =-739;
28248: waveform_sig_rx =-1019;
28249: waveform_sig_rx =-841;
28250: waveform_sig_rx =-919;
28251: waveform_sig_rx =-889;
28252: waveform_sig_rx =-1011;
28253: waveform_sig_rx =-891;
28254: waveform_sig_rx =-850;
28255: waveform_sig_rx =-1159;
28256: waveform_sig_rx =-798;
28257: waveform_sig_rx =-956;
28258: waveform_sig_rx =-1131;
28259: waveform_sig_rx =-832;
28260: waveform_sig_rx =-895;
28261: waveform_sig_rx =-1152;
28262: waveform_sig_rx =-899;
28263: waveform_sig_rx =-868;
28264: waveform_sig_rx =-1180;
28265: waveform_sig_rx =-965;
28266: waveform_sig_rx =-831;
28267: waveform_sig_rx =-1158;
28268: waveform_sig_rx =-1078;
28269: waveform_sig_rx =-791;
28270: waveform_sig_rx =-1132;
28271: waveform_sig_rx =-1082;
28272: waveform_sig_rx =-946;
28273: waveform_sig_rx =-980;
28274: waveform_sig_rx =-1155;
28275: waveform_sig_rx =-952;
28276: waveform_sig_rx =-947;
28277: waveform_sig_rx =-1134;
28278: waveform_sig_rx =-1082;
28279: waveform_sig_rx =-873;
28280: waveform_sig_rx =-1110;
28281: waveform_sig_rx =-1209;
28282: waveform_sig_rx =-823;
28283: waveform_sig_rx =-1096;
28284: waveform_sig_rx =-1230;
28285: waveform_sig_rx =-892;
28286: waveform_sig_rx =-1038;
28287: waveform_sig_rx =-1206;
28288: waveform_sig_rx =-948;
28289: waveform_sig_rx =-1210;
28290: waveform_sig_rx =-962;
28291: waveform_sig_rx =-1133;
28292: waveform_sig_rx =-1036;
28293: waveform_sig_rx =-1177;
28294: waveform_sig_rx =-1050;
28295: waveform_sig_rx =-982;
28296: waveform_sig_rx =-1301;
28297: waveform_sig_rx =-963;
28298: waveform_sig_rx =-1071;
28299: waveform_sig_rx =-1275;
28300: waveform_sig_rx =-972;
28301: waveform_sig_rx =-1020;
28302: waveform_sig_rx =-1320;
28303: waveform_sig_rx =-1004;
28304: waveform_sig_rx =-991;
28305: waveform_sig_rx =-1350;
28306: waveform_sig_rx =-1016;
28307: waveform_sig_rx =-986;
28308: waveform_sig_rx =-1320;
28309: waveform_sig_rx =-1121;
28310: waveform_sig_rx =-975;
28311: waveform_sig_rx =-1239;
28312: waveform_sig_rx =-1156;
28313: waveform_sig_rx =-1112;
28314: waveform_sig_rx =-1024;
28315: waveform_sig_rx =-1285;
28316: waveform_sig_rx =-1061;
28317: waveform_sig_rx =-1014;
28318: waveform_sig_rx =-1292;
28319: waveform_sig_rx =-1164;
28320: waveform_sig_rx =-957;
28321: waveform_sig_rx =-1266;
28322: waveform_sig_rx =-1253;
28323: waveform_sig_rx =-946;
28324: waveform_sig_rx =-1225;
28325: waveform_sig_rx =-1264;
28326: waveform_sig_rx =-1011;
28327: waveform_sig_rx =-1143;
28328: waveform_sig_rx =-1278;
28329: waveform_sig_rx =-1076;
28330: waveform_sig_rx =-1270;
28331: waveform_sig_rx =-1043;
28332: waveform_sig_rx =-1262;
28333: waveform_sig_rx =-1062;
28334: waveform_sig_rx =-1256;
28335: waveform_sig_rx =-1141;
28336: waveform_sig_rx =-1037;
28337: waveform_sig_rx =-1372;
28338: waveform_sig_rx =-1003;
28339: waveform_sig_rx =-1120;
28340: waveform_sig_rx =-1365;
28341: waveform_sig_rx =-981;
28342: waveform_sig_rx =-1084;
28343: waveform_sig_rx =-1430;
28344: waveform_sig_rx =-950;
28345: waveform_sig_rx =-1107;
28346: waveform_sig_rx =-1385;
28347: waveform_sig_rx =-995;
28348: waveform_sig_rx =-1108;
28349: waveform_sig_rx =-1277;
28350: waveform_sig_rx =-1151;
28351: waveform_sig_rx =-1053;
28352: waveform_sig_rx =-1187;
28353: waveform_sig_rx =-1259;
28354: waveform_sig_rx =-1094;
28355: waveform_sig_rx =-1051;
28356: waveform_sig_rx =-1387;
28357: waveform_sig_rx =-1040;
28358: waveform_sig_rx =-1071;
28359: waveform_sig_rx =-1323;
28360: waveform_sig_rx =-1144;
28361: waveform_sig_rx =-984;
28362: waveform_sig_rx =-1271;
28363: waveform_sig_rx =-1235;
28364: waveform_sig_rx =-954;
28365: waveform_sig_rx =-1265;
28366: waveform_sig_rx =-1229;
28367: waveform_sig_rx =-1029;
28368: waveform_sig_rx =-1137;
28369: waveform_sig_rx =-1225;
28370: waveform_sig_rx =-1136;
28371: waveform_sig_rx =-1200;
28372: waveform_sig_rx =-1053;
28373: waveform_sig_rx =-1246;
28374: waveform_sig_rx =-969;
28375: waveform_sig_rx =-1321;
28376: waveform_sig_rx =-1065;
28377: waveform_sig_rx =-1028;
28378: waveform_sig_rx =-1390;
28379: waveform_sig_rx =-887;
28380: waveform_sig_rx =-1163;
28381: waveform_sig_rx =-1323;
28382: waveform_sig_rx =-900;
28383: waveform_sig_rx =-1162;
28384: waveform_sig_rx =-1303;
28385: waveform_sig_rx =-953;
28386: waveform_sig_rx =-1080;
28387: waveform_sig_rx =-1301;
28388: waveform_sig_rx =-1013;
28389: waveform_sig_rx =-1054;
28390: waveform_sig_rx =-1257;
28391: waveform_sig_rx =-1119;
28392: waveform_sig_rx =-997;
28393: waveform_sig_rx =-1167;
28394: waveform_sig_rx =-1219;
28395: waveform_sig_rx =-1008;
28396: waveform_sig_rx =-1016;
28397: waveform_sig_rx =-1331;
28398: waveform_sig_rx =-934;
28399: waveform_sig_rx =-1034;
28400: waveform_sig_rx =-1261;
28401: waveform_sig_rx =-1006;
28402: waveform_sig_rx =-975;
28403: waveform_sig_rx =-1184;
28404: waveform_sig_rx =-1118;
28405: waveform_sig_rx =-919;
28406: waveform_sig_rx =-1108;
28407: waveform_sig_rx =-1188;
28408: waveform_sig_rx =-962;
28409: waveform_sig_rx =-995;
28410: waveform_sig_rx =-1214;
28411: waveform_sig_rx =-987;
28412: waveform_sig_rx =-1090;
28413: waveform_sig_rx =-1022;
28414: waveform_sig_rx =-1099;
28415: waveform_sig_rx =-935;
28416: waveform_sig_rx =-1260;
28417: waveform_sig_rx =-869;
28418: waveform_sig_rx =-1042;
28419: waveform_sig_rx =-1238;
28420: waveform_sig_rx =-787;
28421: waveform_sig_rx =-1137;
28422: waveform_sig_rx =-1129;
28423: waveform_sig_rx =-855;
28424: waveform_sig_rx =-1052;
28425: waveform_sig_rx =-1187;
28426: waveform_sig_rx =-844;
28427: waveform_sig_rx =-984;
28428: waveform_sig_rx =-1175;
28429: waveform_sig_rx =-887;
28430: waveform_sig_rx =-933;
28431: waveform_sig_rx =-1130;
28432: waveform_sig_rx =-1010;
28433: waveform_sig_rx =-848;
28434: waveform_sig_rx =-1046;
28435: waveform_sig_rx =-1101;
28436: waveform_sig_rx =-824;
28437: waveform_sig_rx =-934;
28438: waveform_sig_rx =-1182;
28439: waveform_sig_rx =-738;
28440: waveform_sig_rx =-976;
28441: waveform_sig_rx =-1044;
28442: waveform_sig_rx =-894;
28443: waveform_sig_rx =-869;
28444: waveform_sig_rx =-980;
28445: waveform_sig_rx =-1062;
28446: waveform_sig_rx =-743;
28447: waveform_sig_rx =-952;
28448: waveform_sig_rx =-1099;
28449: waveform_sig_rx =-714;
28450: waveform_sig_rx =-940;
28451: waveform_sig_rx =-1065;
28452: waveform_sig_rx =-768;
28453: waveform_sig_rx =-1020;
28454: waveform_sig_rx =-811;
28455: waveform_sig_rx =-938;
28456: waveform_sig_rx =-811;
28457: waveform_sig_rx =-1038;
28458: waveform_sig_rx =-735;
28459: waveform_sig_rx =-884;
28460: waveform_sig_rx =-1023;
28461: waveform_sig_rx =-663;
28462: waveform_sig_rx =-938;
28463: waveform_sig_rx =-957;
28464: waveform_sig_rx =-655;
28465: waveform_sig_rx =-884;
28466: waveform_sig_rx =-988;
28467: waveform_sig_rx =-678;
28468: waveform_sig_rx =-815;
28469: waveform_sig_rx =-962;
28470: waveform_sig_rx =-744;
28471: waveform_sig_rx =-702;
28472: waveform_sig_rx =-984;
28473: waveform_sig_rx =-818;
28474: waveform_sig_rx =-608;
28475: waveform_sig_rx =-945;
28476: waveform_sig_rx =-816;
28477: waveform_sig_rx =-634;
28478: waveform_sig_rx =-817;
28479: waveform_sig_rx =-867;
28480: waveform_sig_rx =-657;
28481: waveform_sig_rx =-730;
28482: waveform_sig_rx =-857;
28483: waveform_sig_rx =-753;
28484: waveform_sig_rx =-562;
28485: waveform_sig_rx =-863;
28486: waveform_sig_rx =-802;
28487: waveform_sig_rx =-491;
28488: waveform_sig_rx =-822;
28489: waveform_sig_rx =-804;
28490: waveform_sig_rx =-511;
28491: waveform_sig_rx =-736;
28492: waveform_sig_rx =-790;
28493: waveform_sig_rx =-584;
28494: waveform_sig_rx =-816;
28495: waveform_sig_rx =-556;
28496: waveform_sig_rx =-728;
28497: waveform_sig_rx =-586;
28498: waveform_sig_rx =-798;
28499: waveform_sig_rx =-516;
28500: waveform_sig_rx =-651;
28501: waveform_sig_rx =-768;
28502: waveform_sig_rx =-444;
28503: waveform_sig_rx =-688;
28504: waveform_sig_rx =-739;
28505: waveform_sig_rx =-461;
28506: waveform_sig_rx =-613;
28507: waveform_sig_rx =-786;
28508: waveform_sig_rx =-403;
28509: waveform_sig_rx =-572;
28510: waveform_sig_rx =-775;
28511: waveform_sig_rx =-436;
28512: waveform_sig_rx =-473;
28513: waveform_sig_rx =-781;
28514: waveform_sig_rx =-496;
28515: waveform_sig_rx =-413;
28516: waveform_sig_rx =-694;
28517: waveform_sig_rx =-545;
28518: waveform_sig_rx =-476;
28519: waveform_sig_rx =-503;
28520: waveform_sig_rx =-665;
28521: waveform_sig_rx =-431;
28522: waveform_sig_rx =-422;
28523: waveform_sig_rx =-669;
28524: waveform_sig_rx =-459;
28525: waveform_sig_rx =-306;
28526: waveform_sig_rx =-678;
28527: waveform_sig_rx =-474;
28528: waveform_sig_rx =-284;
28529: waveform_sig_rx =-577;
28530: waveform_sig_rx =-514;
28531: waveform_sig_rx =-285;
28532: waveform_sig_rx =-469;
28533: waveform_sig_rx =-524;
28534: waveform_sig_rx =-322;
28535: waveform_sig_rx =-541;
28536: waveform_sig_rx =-294;
28537: waveform_sig_rx =-493;
28538: waveform_sig_rx =-314;
28539: waveform_sig_rx =-542;
28540: waveform_sig_rx =-276;
28541: waveform_sig_rx =-363;
28542: waveform_sig_rx =-530;
28543: waveform_sig_rx =-203;
28544: waveform_sig_rx =-398;
28545: waveform_sig_rx =-534;
28546: waveform_sig_rx =-115;
28547: waveform_sig_rx =-363;
28548: waveform_sig_rx =-550;
28549: waveform_sig_rx =-52;
28550: waveform_sig_rx =-374;
28551: waveform_sig_rx =-457;
28552: waveform_sig_rx =-141;
28553: waveform_sig_rx =-270;
28554: waveform_sig_rx =-441;
28555: waveform_sig_rx =-239;
28556: waveform_sig_rx =-177;
28557: waveform_sig_rx =-357;
28558: waveform_sig_rx =-322;
28559: waveform_sig_rx =-153;
28560: waveform_sig_rx =-213;
28561: waveform_sig_rx =-407;
28562: waveform_sig_rx =-100;
28563: waveform_sig_rx =-152;
28564: waveform_sig_rx =-425;
28565: waveform_sig_rx =-139;
28566: waveform_sig_rx =-53;
28567: waveform_sig_rx =-387;
28568: waveform_sig_rx =-151;
28569: waveform_sig_rx =-49;
28570: waveform_sig_rx =-280;
28571: waveform_sig_rx =-206;
28572: waveform_sig_rx =-33;
28573: waveform_sig_rx =-158;
28574: waveform_sig_rx =-220;
28575: waveform_sig_rx =-77;
28576: waveform_sig_rx =-188;
28577: waveform_sig_rx =-42;
28578: waveform_sig_rx =-193;
28579: waveform_sig_rx =11;
28580: waveform_sig_rx =-303;
28581: waveform_sig_rx =56;
28582: waveform_sig_rx =-100;
28583: waveform_sig_rx =-281;
28584: waveform_sig_rx =161;
28585: waveform_sig_rx =-161;
28586: waveform_sig_rx =-227;
28587: waveform_sig_rx =220;
28588: waveform_sig_rx =-162;
28589: waveform_sig_rx =-227;
28590: waveform_sig_rx =235;
28591: waveform_sig_rx =-145;
28592: waveform_sig_rx =-116;
28593: waveform_sig_rx =103;
28594: waveform_sig_rx =-2;
28595: waveform_sig_rx =-115;
28596: waveform_sig_rx =34;
28597: waveform_sig_rx =121;
28598: waveform_sig_rx =-62;
28599: waveform_sig_rx =-54;
28600: waveform_sig_rx =180;
28601: waveform_sig_rx =37;
28602: waveform_sig_rx =-136;
28603: waveform_sig_rx =244;
28604: waveform_sig_rx =73;
28605: waveform_sig_rx =-117;
28606: waveform_sig_rx =200;
28607: waveform_sig_rx =172;
28608: waveform_sig_rx =-51;
28609: waveform_sig_rx =132;
28610: waveform_sig_rx =224;
28611: waveform_sig_rx =52;
28612: waveform_sig_rx =34;
28613: waveform_sig_rx =266;
28614: waveform_sig_rx =150;
28615: waveform_sig_rx =18;
28616: waveform_sig_rx =234;
28617: waveform_sig_rx =98;
28618: waveform_sig_rx =208;
28619: waveform_sig_rx =118;
28620: waveform_sig_rx =286;
28621: waveform_sig_rx =-5;
28622: waveform_sig_rx =404;
28623: waveform_sig_rx =147;
28624: waveform_sig_rx =30;
28625: waveform_sig_rx =486;
28626: waveform_sig_rx =56;
28627: waveform_sig_rx =125;
28628: waveform_sig_rx =504;
28629: waveform_sig_rx =90;
28630: waveform_sig_rx =162;
28631: waveform_sig_rx =467;
28632: waveform_sig_rx =150;
28633: waveform_sig_rx =215;
28634: waveform_sig_rx =344;
28635: waveform_sig_rx =369;
28636: waveform_sig_rx =119;
28637: waveform_sig_rx =311;
28638: waveform_sig_rx =469;
28639: waveform_sig_rx =163;
28640: waveform_sig_rx =276;
28641: waveform_sig_rx =499;
28642: waveform_sig_rx =284;
28643: waveform_sig_rx =230;
28644: waveform_sig_rx =515;
28645: waveform_sig_rx =333;
28646: waveform_sig_rx =234;
28647: waveform_sig_rx =473;
28648: waveform_sig_rx =459;
28649: waveform_sig_rx =235;
28650: waveform_sig_rx =391;
28651: waveform_sig_rx =511;
28652: waveform_sig_rx =347;
28653: waveform_sig_rx =280;
28654: waveform_sig_rx =590;
28655: waveform_sig_rx =393;
28656: waveform_sig_rx =310;
28657: waveform_sig_rx =553;
28658: waveform_sig_rx =332;
28659: waveform_sig_rx =503;
28660: waveform_sig_rx =450;
28661: waveform_sig_rx =513;
28662: waveform_sig_rx =291;
28663: waveform_sig_rx =694;
28664: waveform_sig_rx =363;
28665: waveform_sig_rx =401;
28666: waveform_sig_rx =720;
28667: waveform_sig_rx =328;
28668: waveform_sig_rx =469;
28669: waveform_sig_rx =694;
28670: waveform_sig_rx =408;
28671: waveform_sig_rx =437;
28672: waveform_sig_rx =715;
28673: waveform_sig_rx =492;
28674: waveform_sig_rx =435;
28675: waveform_sig_rx =631;
28676: waveform_sig_rx =656;
28677: waveform_sig_rx =348;
28678: waveform_sig_rx =659;
28679: waveform_sig_rx =716;
28680: waveform_sig_rx =421;
28681: waveform_sig_rx =600;
28682: waveform_sig_rx =726;
28683: waveform_sig_rx =556;
28684: waveform_sig_rx =505;
28685: waveform_sig_rx =771;
28686: waveform_sig_rx =603;
28687: waveform_sig_rx =491;
28688: waveform_sig_rx =717;
28689: waveform_sig_rx =723;
28690: waveform_sig_rx =505;
28691: waveform_sig_rx =646;
28692: waveform_sig_rx =800;
28693: waveform_sig_rx =569;
28694: waveform_sig_rx =544;
28695: waveform_sig_rx =910;
28696: waveform_sig_rx =570;
28697: waveform_sig_rx =597;
28698: waveform_sig_rx =816;
28699: waveform_sig_rx =524;
28700: waveform_sig_rx =823;
28701: waveform_sig_rx =646;
28702: waveform_sig_rx =739;
28703: waveform_sig_rx =605;
28704: waveform_sig_rx =885;
28705: waveform_sig_rx =625;
28706: waveform_sig_rx =677;
28707: waveform_sig_rx =911;
28708: waveform_sig_rx =642;
28709: waveform_sig_rx =679;
28710: waveform_sig_rx =967;
28711: waveform_sig_rx =665;
28712: waveform_sig_rx =632;
28713: waveform_sig_rx =1001;
28714: waveform_sig_rx =688;
28715: waveform_sig_rx =696;
28716: waveform_sig_rx =907;
28717: waveform_sig_rx =847;
28718: waveform_sig_rx =574;
28719: waveform_sig_rx =925;
28720: waveform_sig_rx =903;
28721: waveform_sig_rx =661;
28722: waveform_sig_rx =842;
28723: waveform_sig_rx =925;
28724: waveform_sig_rx =775;
28725: waveform_sig_rx =742;
28726: waveform_sig_rx =951;
28727: waveform_sig_rx =857;
28728: waveform_sig_rx =707;
28729: waveform_sig_rx =931;
28730: waveform_sig_rx =994;
28731: waveform_sig_rx =650;
28732: waveform_sig_rx =902;
28733: waveform_sig_rx =1047;
28734: waveform_sig_rx =695;
28735: waveform_sig_rx =856;
28736: waveform_sig_rx =1065;
28737: waveform_sig_rx =755;
28738: waveform_sig_rx =909;
28739: waveform_sig_rx =937;
28740: waveform_sig_rx =827;
28741: waveform_sig_rx =1041;
28742: waveform_sig_rx =834;
28743: waveform_sig_rx =1018;
28744: waveform_sig_rx =772;
28745: waveform_sig_rx =1095;
28746: waveform_sig_rx =861;
28747: waveform_sig_rx =839;
28748: waveform_sig_rx =1124;
28749: waveform_sig_rx =805;
28750: waveform_sig_rx =862;
28751: waveform_sig_rx =1190;
28752: waveform_sig_rx =836;
28753: waveform_sig_rx =837;
28754: waveform_sig_rx =1206;
28755: waveform_sig_rx =847;
28756: waveform_sig_rx =844;
28757: waveform_sig_rx =1150;
28758: waveform_sig_rx =964;
28759: waveform_sig_rx =782;
28760: waveform_sig_rx =1130;
28761: waveform_sig_rx =1002;
28762: waveform_sig_rx =903;
28763: waveform_sig_rx =963;
28764: waveform_sig_rx =1091;
28765: waveform_sig_rx =986;
28766: waveform_sig_rx =866;
28767: waveform_sig_rx =1176;
28768: waveform_sig_rx =1010;
28769: waveform_sig_rx =815;
28770: waveform_sig_rx =1170;
28771: waveform_sig_rx =1098;
28772: waveform_sig_rx =800;
28773: waveform_sig_rx =1121;
28774: waveform_sig_rx =1126;
28775: waveform_sig_rx =880;
28776: waveform_sig_rx =1029;
28777: waveform_sig_rx =1170;
28778: waveform_sig_rx =944;
28779: waveform_sig_rx =1037;
28780: waveform_sig_rx =1039;
28781: waveform_sig_rx =1023;
28782: waveform_sig_rx =1100;
28783: waveform_sig_rx =993;
28784: waveform_sig_rx =1149;
28785: waveform_sig_rx =877;
28786: waveform_sig_rx =1281;
28787: waveform_sig_rx =937;
28788: waveform_sig_rx =978;
28789: waveform_sig_rx =1292;
28790: waveform_sig_rx =904;
28791: waveform_sig_rx =1018;
28792: waveform_sig_rx =1331;
28793: waveform_sig_rx =917;
28794: waveform_sig_rx =979;
28795: waveform_sig_rx =1373;
28796: waveform_sig_rx =923;
28797: waveform_sig_rx =1039;
28798: waveform_sig_rx =1286;
28799: waveform_sig_rx =1044;
28800: waveform_sig_rx =974;
28801: waveform_sig_rx =1194;
28802: waveform_sig_rx =1131;
28803: waveform_sig_rx =1052;
28804: waveform_sig_rx =1033;
28805: waveform_sig_rx =1301;
28806: waveform_sig_rx =1020;
28807: waveform_sig_rx =976;
28808: waveform_sig_rx =1346;
28809: waveform_sig_rx =1019;
28810: waveform_sig_rx =1004;
28811: waveform_sig_rx =1260;
28812: waveform_sig_rx =1148;
28813: waveform_sig_rx =961;
28814: waveform_sig_rx =1182;
28815: waveform_sig_rx =1234;
28816: waveform_sig_rx =994;
28817: waveform_sig_rx =1118;
28818: waveform_sig_rx =1280;
28819: waveform_sig_rx =1032;
28820: waveform_sig_rx =1116;
28821: waveform_sig_rx =1110;
28822: waveform_sig_rx =1132;
28823: waveform_sig_rx =1145;
28824: waveform_sig_rx =1114;
28825: waveform_sig_rx =1212;
28826: waveform_sig_rx =937;
28827: waveform_sig_rx =1409;
28828: waveform_sig_rx =957;
28829: waveform_sig_rx =1098;
28830: waveform_sig_rx =1383;
28831: waveform_sig_rx =890;
28832: waveform_sig_rx =1173;
28833: waveform_sig_rx =1337;
28834: waveform_sig_rx =955;
28835: waveform_sig_rx =1135;
28836: waveform_sig_rx =1318;
28837: waveform_sig_rx =1004;
28838: waveform_sig_rx =1097;
28839: waveform_sig_rx =1260;
28840: waveform_sig_rx =1124;
28841: waveform_sig_rx =994;
28842: waveform_sig_rx =1257;
28843: waveform_sig_rx =1209;
28844: waveform_sig_rx =1041;
28845: waveform_sig_rx =1101;
28846: waveform_sig_rx =1333;
28847: waveform_sig_rx =1014;
28848: waveform_sig_rx =1060;
28849: waveform_sig_rx =1368;
28850: waveform_sig_rx =1023;
28851: waveform_sig_rx =1076;
28852: waveform_sig_rx =1280;
28853: waveform_sig_rx =1149;
28854: waveform_sig_rx =1034;
28855: waveform_sig_rx =1182;
28856: waveform_sig_rx =1266;
28857: waveform_sig_rx =1040;
28858: waveform_sig_rx =1082;
28859: waveform_sig_rx =1331;
28860: waveform_sig_rx =1029;
28861: waveform_sig_rx =1118;
28862: waveform_sig_rx =1197;
28863: waveform_sig_rx =1108;
28864: waveform_sig_rx =1173;
28865: waveform_sig_rx =1171;
28866: waveform_sig_rx =1129;
28867: waveform_sig_rx =1011;
28868: waveform_sig_rx =1398;
28869: waveform_sig_rx =890;
28870: waveform_sig_rx =1178;
28871: waveform_sig_rx =1287;
28872: waveform_sig_rx =914;
28873: waveform_sig_rx =1200;
28874: waveform_sig_rx =1263;
28875: waveform_sig_rx =988;
28876: waveform_sig_rx =1081;
28877: waveform_sig_rx =1312;
28878: waveform_sig_rx =996;
28879: waveform_sig_rx =1063;
28880: waveform_sig_rx =1246;
28881: waveform_sig_rx =1105;
28882: waveform_sig_rx =952;
28883: waveform_sig_rx =1248;
28884: waveform_sig_rx =1153;
28885: waveform_sig_rx =975;
28886: waveform_sig_rx =1101;
28887: waveform_sig_rx =1292;
28888: waveform_sig_rx =948;
28889: waveform_sig_rx =1088;
28890: waveform_sig_rx =1276;
28891: waveform_sig_rx =988;
28892: waveform_sig_rx =1077;
28893: waveform_sig_rx =1180;
28894: waveform_sig_rx =1153;
28895: waveform_sig_rx =960;
28896: waveform_sig_rx =1104;
28897: waveform_sig_rx =1267;
28898: waveform_sig_rx =889;
28899: waveform_sig_rx =1089;
28900: waveform_sig_rx =1320;
28901: waveform_sig_rx =870;
28902: waveform_sig_rx =1146;
28903: waveform_sig_rx =1057;
28904: waveform_sig_rx =1013;
28905: waveform_sig_rx =1143;
28906: waveform_sig_rx =1032;
28907: waveform_sig_rx =1071;
28908: waveform_sig_rx =969;
28909: waveform_sig_rx =1253;
28910: waveform_sig_rx =842;
28911: waveform_sig_rx =1075;
28912: waveform_sig_rx =1177;
28913: waveform_sig_rx =875;
28914: waveform_sig_rx =1081;
28915: waveform_sig_rx =1175;
28916: waveform_sig_rx =897;
28917: waveform_sig_rx =992;
28918: waveform_sig_rx =1231;
28919: waveform_sig_rx =916;
28920: waveform_sig_rx =960;
28921: waveform_sig_rx =1193;
28922: waveform_sig_rx =1012;
28923: waveform_sig_rx =808;
28924: waveform_sig_rx =1207;
28925: waveform_sig_rx =1007;
28926: waveform_sig_rx =871;
28927: waveform_sig_rx =1074;
28928: waveform_sig_rx =1094;
28929: waveform_sig_rx =872;
28930: waveform_sig_rx =991;
28931: waveform_sig_rx =1090;
28932: waveform_sig_rx =955;
28933: waveform_sig_rx =858;
28934: waveform_sig_rx =1074;
28935: waveform_sig_rx =1080;
28936: waveform_sig_rx =735;
28937: waveform_sig_rx =1087;
28938: waveform_sig_rx =1078;
28939: waveform_sig_rx =732;
28940: waveform_sig_rx =1028;
28941: waveform_sig_rx =1069;
28942: waveform_sig_rx =799;
28943: waveform_sig_rx =1035;
28944: waveform_sig_rx =887;
28945: waveform_sig_rx =931;
28946: waveform_sig_rx =965;
28947: waveform_sig_rx =894;
28948: waveform_sig_rx =950;
28949: waveform_sig_rx =817;
28950: waveform_sig_rx =1110;
28951: waveform_sig_rx =724;
28952: waveform_sig_rx =939;
28953: waveform_sig_rx =1014;
28954: waveform_sig_rx =750;
28955: waveform_sig_rx =897;
28956: waveform_sig_rx =1034;
28957: waveform_sig_rx =729;
28958: waveform_sig_rx =783;
28959: waveform_sig_rx =1107;
28960: waveform_sig_rx =668;
28961: waveform_sig_rx =797;
28962: waveform_sig_rx =1078;
28963: waveform_sig_rx =731;
28964: waveform_sig_rx =716;
28965: waveform_sig_rx =1028;
28966: waveform_sig_rx =766;
28967: waveform_sig_rx =769;
28968: waveform_sig_rx =811;
28969: waveform_sig_rx =940;
28970: waveform_sig_rx =717;
28971: waveform_sig_rx =756;
28972: waveform_sig_rx =973;
28973: waveform_sig_rx =737;
28974: waveform_sig_rx =661;
28975: waveform_sig_rx =951;
28976: waveform_sig_rx =805;
28977: waveform_sig_rx =577;
28978: waveform_sig_rx =930;
28979: waveform_sig_rx =814;
28980: waveform_sig_rx =585;
28981: waveform_sig_rx =836;
28982: waveform_sig_rx =846;
28983: waveform_sig_rx =605;
28984: waveform_sig_rx =795;
28985: waveform_sig_rx =661;
28986: waveform_sig_rx =771;
28987: waveform_sig_rx =727;
28988: waveform_sig_rx =706;
28989: waveform_sig_rx =747;
28990: waveform_sig_rx =568;
28991: waveform_sig_rx =895;
28992: waveform_sig_rx =527;
28993: waveform_sig_rx =680;
28994: waveform_sig_rx =855;
28995: waveform_sig_rx =491;
28996: waveform_sig_rx =668;
28997: waveform_sig_rx =885;
28998: waveform_sig_rx =427;
28999: waveform_sig_rx =642;
29000: waveform_sig_rx =896;
29001: waveform_sig_rx =390;
29002: waveform_sig_rx =687;
29003: waveform_sig_rx =784;
29004: waveform_sig_rx =517;
29005: waveform_sig_rx =573;
29006: waveform_sig_rx =730;
29007: waveform_sig_rx =577;
29008: waveform_sig_rx =548;
29009: waveform_sig_rx =557;
29010: waveform_sig_rx =776;
29011: waveform_sig_rx =421;
29012: waveform_sig_rx =540;
29013: waveform_sig_rx =757;
29014: waveform_sig_rx =425;
29015: waveform_sig_rx =469;
29016: waveform_sig_rx =720;
29017: waveform_sig_rx =527;
29018: waveform_sig_rx =380;
29019: waveform_sig_rx =679;
29020: waveform_sig_rx =528;
29021: waveform_sig_rx =375;
29022: waveform_sig_rx =561;
29023: waveform_sig_rx =610;
29024: waveform_sig_rx =393;
29025: waveform_sig_rx =534;
29026: waveform_sig_rx =447;
29027: waveform_sig_rx =525;
29028: waveform_sig_rx =430;
29029: waveform_sig_rx =504;
29030: waveform_sig_rx =452;
29031: waveform_sig_rx =309;
29032: waveform_sig_rx =701;
29033: waveform_sig_rx =201;
29034: waveform_sig_rx =480;
29035: waveform_sig_rx =603;
29036: waveform_sig_rx =141;
29037: waveform_sig_rx =518;
29038: waveform_sig_rx =579;
29039: waveform_sig_rx =128;
29040: waveform_sig_rx =476;
29041: waveform_sig_rx =543;
29042: waveform_sig_rx =157;
29043: waveform_sig_rx =425;
29044: waveform_sig_rx =447;
29045: waveform_sig_rx =302;
29046: waveform_sig_rx =233;
29047: waveform_sig_rx =470;
29048: waveform_sig_rx =345;
29049: waveform_sig_rx =211;
29050: waveform_sig_rx =312;
29051: waveform_sig_rx =460;
29052: waveform_sig_rx =97;
29053: waveform_sig_rx =290;
29054: waveform_sig_rx =461;
29055: waveform_sig_rx =117;
29056: waveform_sig_rx =213;
29057: waveform_sig_rx =409;
29058: waveform_sig_rx =198;
29059: waveform_sig_rx =138;
29060: waveform_sig_rx =340;
29061: waveform_sig_rx =265;
29062: waveform_sig_rx =111;
29063: waveform_sig_rx =213;
29064: waveform_sig_rx =382;
29065: waveform_sig_rx =57;
29066: waveform_sig_rx =228;
29067: waveform_sig_rx =203;
29068: waveform_sig_rx =179;
29069: waveform_sig_rx =166;
29070: waveform_sig_rx =225;
29071: waveform_sig_rx =93;
29072: waveform_sig_rx =103;
29073: waveform_sig_rx =380;
29074: waveform_sig_rx =-138;
29075: waveform_sig_rx =252;
29076: waveform_sig_rx =262;
29077: waveform_sig_rx =-144;
29078: waveform_sig_rx =258;
29079: waveform_sig_rx =211;
29080: waveform_sig_rx =-144;
29081: waveform_sig_rx =203;
29082: waveform_sig_rx =165;
29083: waveform_sig_rx =-73;
29084: waveform_sig_rx =83;
29085: waveform_sig_rx =125;
29086: waveform_sig_rx =38;
29087: waveform_sig_rx =-148;
29088: waveform_sig_rx =225;
29089: waveform_sig_rx =33;
29090: waveform_sig_rx =-144;
29091: waveform_sig_rx =107;
29092: waveform_sig_rx =120;
29093: waveform_sig_rx =-177;
29094: waveform_sig_rx =53;
29095: waveform_sig_rx =112;
29096: waveform_sig_rx =-149;
29097: waveform_sig_rx =-76;
29098: waveform_sig_rx =112;
29099: waveform_sig_rx =-82;
29100: waveform_sig_rx =-174;
29101: waveform_sig_rx =32;
29102: waveform_sig_rx =-21;
29103: waveform_sig_rx =-227;
29104: waveform_sig_rx =-77;
29105: waveform_sig_rx =115;
29106: waveform_sig_rx =-337;
29107: waveform_sig_rx =-41;
29108: waveform_sig_rx =-134;
29109: waveform_sig_rx =-173;
29110: waveform_sig_rx =-78;
29111: waveform_sig_rx =-111;
29112: waveform_sig_rx =-241;
29113: waveform_sig_rx =-139;
29114: waveform_sig_rx =-13;
29115: waveform_sig_rx =-400;
29116: waveform_sig_rx =-31;
29117: waveform_sig_rx =-141;
29118: waveform_sig_rx =-368;
29119: waveform_sig_rx =-82;
29120: waveform_sig_rx =-113;
29121: waveform_sig_rx =-383;
29122: waveform_sig_rx =-175;
29123: waveform_sig_rx =-95;
29124: waveform_sig_rx =-395;
29125: waveform_sig_rx =-244;
29126: waveform_sig_rx =-112;
29127: waveform_sig_rx =-331;
29128: waveform_sig_rx =-445;
29129: waveform_sig_rx =-43;
29130: waveform_sig_rx =-360;
29131: waveform_sig_rx =-397;
29132: waveform_sig_rx =-209;
29133: waveform_sig_rx =-245;
29134: waveform_sig_rx =-468;
29135: waveform_sig_rx =-286;
29136: waveform_sig_rx =-221;
29137: waveform_sig_rx =-417;
29138: waveform_sig_rx =-396;
29139: waveform_sig_rx =-214;
29140: waveform_sig_rx =-370;
29141: waveform_sig_rx =-525;
29142: waveform_sig_rx =-237;
29143: waveform_sig_rx =-316;
29144: waveform_sig_rx =-576;
29145: waveform_sig_rx =-310;
29146: waveform_sig_rx =-243;
29147: waveform_sig_rx =-641;
29148: waveform_sig_rx =-255;
29149: waveform_sig_rx =-499;
29150: waveform_sig_rx =-435;
29151: waveform_sig_rx =-383;
29152: waveform_sig_rx =-476;
29153: waveform_sig_rx =-479;
29154: waveform_sig_rx =-471;
29155: waveform_sig_rx =-365;
29156: waveform_sig_rx =-617;
29157: waveform_sig_rx =-411;
29158: waveform_sig_rx =-401;
29159: waveform_sig_rx =-657;
29160: waveform_sig_rx =-432;
29161: waveform_sig_rx =-334;
29162: waveform_sig_rx =-757;
29163: waveform_sig_rx =-435;
29164: waveform_sig_rx =-369;
29165: waveform_sig_rx =-752;
29166: waveform_sig_rx =-485;
29167: waveform_sig_rx =-424;
29168: waveform_sig_rx =-639;
29169: waveform_sig_rx =-687;
29170: waveform_sig_rx =-347;
29171: waveform_sig_rx =-642;
29172: waveform_sig_rx =-691;
29173: waveform_sig_rx =-495;
29174: waveform_sig_rx =-545;
29175: waveform_sig_rx =-719;
29176: waveform_sig_rx =-582;
29177: waveform_sig_rx =-504;
29178: waveform_sig_rx =-676;
29179: waveform_sig_rx =-750;
29180: waveform_sig_rx =-420;
29181: waveform_sig_rx =-665;
29182: waveform_sig_rx =-852;
29183: waveform_sig_rx =-403;
29184: waveform_sig_rx =-662;
29185: waveform_sig_rx =-840;
29186: waveform_sig_rx =-519;
29187: waveform_sig_rx =-617;
29188: waveform_sig_rx =-795;
29189: waveform_sig_rx =-567;
29190: waveform_sig_rx =-810;
29191: waveform_sig_rx =-600;
29192: waveform_sig_rx =-741;
29193: waveform_sig_rx =-668;
29194: waveform_sig_rx =-724;
29195: waveform_sig_rx =-777;
29196: waveform_sig_rx =-541;
29197: waveform_sig_rx =-943;
29198: waveform_sig_rx =-678;
29199: waveform_sig_rx =-614;
29200: waveform_sig_rx =-981;
29201: waveform_sig_rx =-631;
29202: waveform_sig_rx =-626;
29203: waveform_sig_rx =-1021;
29204: waveform_sig_rx =-670;
29205: waveform_sig_rx =-627;
29206: waveform_sig_rx =-998;
29207: waveform_sig_rx =-726;
29208: waveform_sig_rx =-645;
29209: waveform_sig_rx =-921;
29210: waveform_sig_rx =-879;
29211: waveform_sig_rx =-623;
29212: waveform_sig_rx =-915;
29213: waveform_sig_rx =-866;
29214: waveform_sig_rx =-809;
29215: waveform_sig_rx =-729;
29216: waveform_sig_rx =-957;
29217: waveform_sig_rx =-872;
29218: waveform_sig_rx =-655;
29219: waveform_sig_rx =-1011;
29220: waveform_sig_rx =-936;
29221: waveform_sig_rx =-618;
29222: waveform_sig_rx =-994;
29223: waveform_sig_rx =-955;
29224: waveform_sig_rx =-705;
29225: waveform_sig_rx =-929;
29226: waveform_sig_rx =-992;
29227: waveform_sig_rx =-838;
29228: waveform_sig_rx =-801;
29229: waveform_sig_rx =-1042;
29230: waveform_sig_rx =-839;
29231: waveform_sig_rx =-981;
29232: waveform_sig_rx =-845;
29233: waveform_sig_rx =-982;
29234: waveform_sig_rx =-848;
29235: waveform_sig_rx =-1008;
29236: waveform_sig_rx =-967;
29237: waveform_sig_rx =-763;
29238: waveform_sig_rx =-1174;
29239: waveform_sig_rx =-804;
29240: waveform_sig_rx =-825;
29241: waveform_sig_rx =-1199;
29242: waveform_sig_rx =-787;
29243: waveform_sig_rx =-843;
29244: waveform_sig_rx =-1251;
29245: waveform_sig_rx =-810;
29246: waveform_sig_rx =-878;
29247: waveform_sig_rx =-1217;
29248: waveform_sig_rx =-863;
29249: waveform_sig_rx =-912;
29250: waveform_sig_rx =-1112;
29251: waveform_sig_rx =-1039;
29252: waveform_sig_rx =-872;
29253: waveform_sig_rx =-1029;
29254: waveform_sig_rx =-1090;
29255: waveform_sig_rx =-1003;
29256: waveform_sig_rx =-839;
29257: waveform_sig_rx =-1247;
29258: waveform_sig_rx =-968;
29259: waveform_sig_rx =-872;
29260: waveform_sig_rx =-1250;
29261: waveform_sig_rx =-1010;
29262: waveform_sig_rx =-896;
29263: waveform_sig_rx =-1155;
29264: waveform_sig_rx =-1127;
29265: waveform_sig_rx =-954;
29266: waveform_sig_rx =-1031;
29267: waveform_sig_rx =-1207;
29268: waveform_sig_rx =-989;
29269: waveform_sig_rx =-951;
29270: waveform_sig_rx =-1231;
29271: waveform_sig_rx =-964;
29272: waveform_sig_rx =-1147;
29273: waveform_sig_rx =-1000;
29274: waveform_sig_rx =-1144;
29275: waveform_sig_rx =-988;
29276: waveform_sig_rx =-1201;
29277: waveform_sig_rx =-1078;
29278: waveform_sig_rx =-931;
29279: waveform_sig_rx =-1356;
29280: waveform_sig_rx =-932;
29281: waveform_sig_rx =-1027;
29282: waveform_sig_rx =-1367;
29283: waveform_sig_rx =-875;
29284: waveform_sig_rx =-1074;
29285: waveform_sig_rx =-1331;
29286: waveform_sig_rx =-915;
29287: waveform_sig_rx =-1090;
29288: waveform_sig_rx =-1249;
29289: waveform_sig_rx =-1041;
29290: waveform_sig_rx =-1044;
29291: waveform_sig_rx =-1185;
29292: waveform_sig_rx =-1244;
29293: waveform_sig_rx =-938;
29294: waveform_sig_rx =-1177;
29295: waveform_sig_rx =-1281;
29296: waveform_sig_rx =-1038;
29297: waveform_sig_rx =-1070;
29298: waveform_sig_rx =-1357;
29299: waveform_sig_rx =-1039;
29300: waveform_sig_rx =-1064;
29301: waveform_sig_rx =-1301;
29302: waveform_sig_rx =-1131;
29303: waveform_sig_rx =-1016;
29304: waveform_sig_rx =-1222;
29305: waveform_sig_rx =-1258;
29306: waveform_sig_rx =-1017;
29307: waveform_sig_rx =-1143;
29308: waveform_sig_rx =-1302;
29309: waveform_sig_rx =-1050;
29310: waveform_sig_rx =-1036;
29311: waveform_sig_rx =-1328;
29312: waveform_sig_rx =-1033;
29313: waveform_sig_rx =-1221;
29314: waveform_sig_rx =-1111;
29315: waveform_sig_rx =-1177;
29316: waveform_sig_rx =-1055;
29317: waveform_sig_rx =-1313;
29318: waveform_sig_rx =-1070;
29319: waveform_sig_rx =-1052;
29320: waveform_sig_rx =-1412;
29321: waveform_sig_rx =-938;
29322: waveform_sig_rx =-1198;
29323: waveform_sig_rx =-1331;
29324: waveform_sig_rx =-981;
29325: waveform_sig_rx =-1160;
29326: waveform_sig_rx =-1316;
29327: waveform_sig_rx =-1046;
29328: waveform_sig_rx =-1090;
29329: waveform_sig_rx =-1323;
29330: waveform_sig_rx =-1118;
29331: waveform_sig_rx =-1032;
29332: waveform_sig_rx =-1303;
29333: waveform_sig_rx =-1234;
29334: waveform_sig_rx =-969;
29335: waveform_sig_rx =-1272;
29336: waveform_sig_rx =-1253;
29337: waveform_sig_rx =-1034;
29338: waveform_sig_rx =-1086;
29339: waveform_sig_rx =-1346;
29340: waveform_sig_rx =-1012;
29341: waveform_sig_rx =-1110;
29342: waveform_sig_rx =-1271;
29343: waveform_sig_rx =-1141;
29344: waveform_sig_rx =-1053;
29345: waveform_sig_rx =-1181;
29346: waveform_sig_rx =-1293;
29347: waveform_sig_rx =-970;
29348: waveform_sig_rx =-1147;
29349: waveform_sig_rx =-1351;
29350: waveform_sig_rx =-971;
29351: waveform_sig_rx =-1088;
29352: waveform_sig_rx =-1307;
29353: waveform_sig_rx =-995;
29354: waveform_sig_rx =-1266;
29355: waveform_sig_rx =-1075;
29356: waveform_sig_rx =-1180;
29357: waveform_sig_rx =-1079;
29358: waveform_sig_rx =-1266;
29359: waveform_sig_rx =-1054;
29360: waveform_sig_rx =-1086;
29361: waveform_sig_rx =-1328;
29362: waveform_sig_rx =-968;
29363: waveform_sig_rx =-1181;
29364: waveform_sig_rx =-1269;
29365: waveform_sig_rx =-995;
29366: waveform_sig_rx =-1089;
29367: waveform_sig_rx =-1310;
29368: waveform_sig_rx =-1004;
29369: waveform_sig_rx =-1017;
29370: waveform_sig_rx =-1313;
29371: waveform_sig_rx =-1017;
29372: waveform_sig_rx =-977;
29373: waveform_sig_rx =-1293;
29374: waveform_sig_rx =-1114;
29375: waveform_sig_rx =-933;
29376: waveform_sig_rx =-1216;
29377: waveform_sig_rx =-1154;
29378: waveform_sig_rx =-998;
29379: waveform_sig_rx =-1051;
29380: waveform_sig_rx =-1254;
29381: waveform_sig_rx =-987;
29382: waveform_sig_rx =-1034;
29383: waveform_sig_rx =-1188;
29384: waveform_sig_rx =-1096;
29385: waveform_sig_rx =-927;
29386: waveform_sig_rx =-1144;
29387: waveform_sig_rx =-1236;
29388: waveform_sig_rx =-831;
29389: waveform_sig_rx =-1160;
29390: waveform_sig_rx =-1238;
29391: waveform_sig_rx =-864;
29392: waveform_sig_rx =-1102;
29393: waveform_sig_rx =-1153;
29394: waveform_sig_rx =-954;
29395: waveform_sig_rx =-1214;
29396: waveform_sig_rx =-928;
29397: waveform_sig_rx =-1141;
29398: waveform_sig_rx =-947;
29399: waveform_sig_rx =-1170;
29400: waveform_sig_rx =-990;
29401: waveform_sig_rx =-966;
29402: waveform_sig_rx =-1241;
29403: waveform_sig_rx =-874;
29404: waveform_sig_rx =-1033;
29405: waveform_sig_rx =-1192;
29406: waveform_sig_rx =-861;
29407: waveform_sig_rx =-962;
29408: waveform_sig_rx =-1234;
29409: waveform_sig_rx =-865;
29410: waveform_sig_rx =-915;
29411: waveform_sig_rx =-1236;
29412: waveform_sig_rx =-864;
29413: waveform_sig_rx =-896;
29414: waveform_sig_rx =-1189;
29415: waveform_sig_rx =-934;
29416: waveform_sig_rx =-863;
29417: waveform_sig_rx =-1053;
29418: waveform_sig_rx =-1010;
29419: waveform_sig_rx =-928;
29420: waveform_sig_rx =-871;
29421: waveform_sig_rx =-1164;
29422: waveform_sig_rx =-848;
29423: waveform_sig_rx =-862;
29424: waveform_sig_rx =-1117;
29425: waveform_sig_rx =-903;
29426: waveform_sig_rx =-778;
29427: waveform_sig_rx =-1073;
29428: waveform_sig_rx =-1030;
29429: waveform_sig_rx =-728;
29430: waveform_sig_rx =-1029;
29431: waveform_sig_rx =-1027;
29432: waveform_sig_rx =-750;
29433: waveform_sig_rx =-964;
29434: waveform_sig_rx =-996;
29435: waveform_sig_rx =-838;
29436: waveform_sig_rx =-1015;
29437: waveform_sig_rx =-763;
29438: waveform_sig_rx =-1015;
29439: waveform_sig_rx =-748;
29440: waveform_sig_rx =-1039;
29441: waveform_sig_rx =-835;
29442: waveform_sig_rx =-775;
29443: waveform_sig_rx =-1100;
29444: waveform_sig_rx =-665;
29445: waveform_sig_rx =-840;
29446: waveform_sig_rx =-1072;
29447: waveform_sig_rx =-613;
29448: waveform_sig_rx =-838;
29449: waveform_sig_rx =-1062;
29450: waveform_sig_rx =-616;
29451: waveform_sig_rx =-813;
29452: waveform_sig_rx =-1006;
29453: waveform_sig_rx =-673;
29454: waveform_sig_rx =-776;
29455: waveform_sig_rx =-956;
29456: waveform_sig_rx =-755;
29457: waveform_sig_rx =-704;
29458: waveform_sig_rx =-871;
29459: waveform_sig_rx =-868;
29460: waveform_sig_rx =-717;
29461: waveform_sig_rx =-685;
29462: waveform_sig_rx =-1000;
29463: waveform_sig_rx =-615;
29464: waveform_sig_rx =-698;
29465: waveform_sig_rx =-962;
29466: waveform_sig_rx =-690;
29467: waveform_sig_rx =-625;
29468: waveform_sig_rx =-884;
29469: waveform_sig_rx =-761;
29470: waveform_sig_rx =-589;
29471: waveform_sig_rx =-780;
29472: waveform_sig_rx =-790;
29473: waveform_sig_rx =-584;
29474: waveform_sig_rx =-650;
29475: waveform_sig_rx =-787;
29476: waveform_sig_rx =-617;
29477: waveform_sig_rx =-727;
29478: waveform_sig_rx =-597;
29479: waveform_sig_rx =-766;
29480: waveform_sig_rx =-505;
29481: waveform_sig_rx =-874;
29482: waveform_sig_rx =-516;
29483: waveform_sig_rx =-602;
29484: waveform_sig_rx =-889;
29485: waveform_sig_rx =-386;
29486: waveform_sig_rx =-709;
29487: waveform_sig_rx =-810;
29488: waveform_sig_rx =-376;
29489: waveform_sig_rx =-683;
29490: waveform_sig_rx =-773;
29491: waveform_sig_rx =-389;
29492: waveform_sig_rx =-629;
29493: waveform_sig_rx =-710;
29494: waveform_sig_rx =-473;
29495: waveform_sig_rx =-530;
29496: waveform_sig_rx =-689;
29497: waveform_sig_rx =-571;
29498: waveform_sig_rx =-420;
29499: waveform_sig_rx =-612;
29500: waveform_sig_rx =-663;
29501: waveform_sig_rx =-402;
29502: waveform_sig_rx =-500;
29503: waveform_sig_rx =-747;
29504: waveform_sig_rx =-308;
29505: waveform_sig_rx =-503;
29506: waveform_sig_rx =-651;
29507: waveform_sig_rx =-410;
29508: waveform_sig_rx =-409;
29509: waveform_sig_rx =-582;
29510: waveform_sig_rx =-513;
29511: waveform_sig_rx =-339;
29512: waveform_sig_rx =-498;
29513: waveform_sig_rx =-584;
29514: waveform_sig_rx =-298;
29515: waveform_sig_rx =-388;
29516: waveform_sig_rx =-589;
29517: waveform_sig_rx =-316;
29518: waveform_sig_rx =-499;
29519: waveform_sig_rx =-369;
29520: waveform_sig_rx =-430;
29521: waveform_sig_rx =-306;
29522: waveform_sig_rx =-585;
29523: waveform_sig_rx =-198;
29524: waveform_sig_rx =-419;
29525: waveform_sig_rx =-552;
29526: waveform_sig_rx =-121;
29527: waveform_sig_rx =-488;
29528: waveform_sig_rx =-454;
29529: waveform_sig_rx =-116;
29530: waveform_sig_rx =-426;
29531: waveform_sig_rx =-470;
29532: waveform_sig_rx =-137;
29533: waveform_sig_rx =-361;
29534: waveform_sig_rx =-414;
29535: waveform_sig_rx =-229;
29536: waveform_sig_rx =-228;
29537: waveform_sig_rx =-433;
29538: waveform_sig_rx =-331;
29539: waveform_sig_rx =-90;
29540: waveform_sig_rx =-413;
29541: waveform_sig_rx =-359;
29542: waveform_sig_rx =-80;
29543: waveform_sig_rx =-315;
29544: waveform_sig_rx =-393;
29545: waveform_sig_rx =-65;
29546: waveform_sig_rx =-262;
29547: waveform_sig_rx =-321;
29548: waveform_sig_rx =-184;
29549: waveform_sig_rx =-92;
29550: waveform_sig_rx =-300;
29551: waveform_sig_rx =-273;
29552: waveform_sig_rx =0;
29553: waveform_sig_rx =-260;
29554: waveform_sig_rx =-300;
29555: waveform_sig_rx =25;
29556: waveform_sig_rx =-184;
29557: waveform_sig_rx =-275;
29558: waveform_sig_rx =-9;
29559: waveform_sig_rx =-245;
29560: waveform_sig_rx =-56;
29561: waveform_sig_rx =-132;
29562: waveform_sig_rx =-54;
29563: waveform_sig_rx =-256;
29564: waveform_sig_rx =87;
29565: waveform_sig_rx =-173;
29566: waveform_sig_rx =-189;
29567: waveform_sig_rx =121;
29568: waveform_sig_rx =-197;
29569: waveform_sig_rx =-125;
29570: waveform_sig_rx =93;
29571: waveform_sig_rx =-86;
29572: waveform_sig_rx =-189;
29573: waveform_sig_rx =136;
29574: waveform_sig_rx =-23;
29575: waveform_sig_rx =-164;
29576: waveform_sig_rx =94;
29577: waveform_sig_rx =81;
29578: waveform_sig_rx =-209;
29579: waveform_sig_rx =49;
29580: waveform_sig_rx =172;
29581: waveform_sig_rx =-137;
29582: waveform_sig_rx =24;
29583: waveform_sig_rx =160;
29584: waveform_sig_rx =6;
29585: waveform_sig_rx =-66;
29586: waveform_sig_rx =163;
29587: waveform_sig_rx =74;
29588: waveform_sig_rx =-51;
29589: waveform_sig_rx =105;
29590: waveform_sig_rx =231;
29591: waveform_sig_rx =-44;
29592: waveform_sig_rx =53;
29593: waveform_sig_rx =306;
29594: waveform_sig_rx =5;
29595: waveform_sig_rx =9;
29596: waveform_sig_rx =335;
29597: waveform_sig_rx =68;
29598: waveform_sig_rx =64;
29599: waveform_sig_rx =274;
29600: waveform_sig_rx =-1;
29601: waveform_sig_rx =301;
29602: waveform_sig_rx =110;
29603: waveform_sig_rx =223;
29604: waveform_sig_rx =79;
29605: waveform_sig_rx =321;
29606: waveform_sig_rx =160;
29607: waveform_sig_rx =113;
29608: waveform_sig_rx =361;
29609: waveform_sig_rx =181;
29610: waveform_sig_rx =91;
29611: waveform_sig_rx =423;
29612: waveform_sig_rx =215;
29613: waveform_sig_rx =25;
29614: waveform_sig_rx =513;
29615: waveform_sig_rx =205;
29616: waveform_sig_rx =109;
29617: waveform_sig_rx =431;
29618: waveform_sig_rx =325;
29619: waveform_sig_rx =108;
29620: waveform_sig_rx =371;
29621: waveform_sig_rx =422;
29622: waveform_sig_rx =188;
29623: waveform_sig_rx =308;
29624: waveform_sig_rx =437;
29625: waveform_sig_rx =320;
29626: waveform_sig_rx =243;
29627: waveform_sig_rx =465;
29628: waveform_sig_rx =401;
29629: waveform_sig_rx =224;
29630: waveform_sig_rx =410;
29631: waveform_sig_rx =574;
29632: waveform_sig_rx =197;
29633: waveform_sig_rx =401;
29634: waveform_sig_rx =596;
29635: waveform_sig_rx =236;
29636: waveform_sig_rx =357;
29637: waveform_sig_rx =578;
29638: waveform_sig_rx =334;
29639: waveform_sig_rx =393;
29640: waveform_sig_rx =468;
29641: waveform_sig_rx =343;
29642: waveform_sig_rx =574;
29643: waveform_sig_rx =332;
29644: waveform_sig_rx =588;
29645: waveform_sig_rx =314;
29646: waveform_sig_rx =589;
29647: waveform_sig_rx =496;
29648: waveform_sig_rx =313;
29649: waveform_sig_rx =718;
29650: waveform_sig_rx =428;
29651: waveform_sig_rx =327;
29652: waveform_sig_rx =795;
29653: waveform_sig_rx =404;
29654: waveform_sig_rx =353;
29655: waveform_sig_rx =806;
29656: waveform_sig_rx =421;
29657: waveform_sig_rx =434;
29658: waveform_sig_rx =683;
29659: waveform_sig_rx =596;
29660: waveform_sig_rx =389;
29661: waveform_sig_rx =651;
29662: waveform_sig_rx =657;
29663: waveform_sig_rx =455;
29664: waveform_sig_rx =577;
29665: waveform_sig_rx =686;
29666: waveform_sig_rx =610;
29667: waveform_sig_rx =471;
29668: waveform_sig_rx =752;
29669: waveform_sig_rx =715;
29670: waveform_sig_rx =399;
29671: waveform_sig_rx =768;
29672: waveform_sig_rx =781;
29673: waveform_sig_rx =401;
29674: waveform_sig_rx =754;
29675: waveform_sig_rx =753;
29676: waveform_sig_rx =551;
29677: waveform_sig_rx =648;
29678: waveform_sig_rx =783;
29679: waveform_sig_rx =678;
29680: waveform_sig_rx =587;
29681: waveform_sig_rx =740;
29682: waveform_sig_rx =645;
29683: waveform_sig_rx =733;
29684: waveform_sig_rx =643;
29685: waveform_sig_rx =793;
29686: waveform_sig_rx =504;
29687: waveform_sig_rx =926;
29688: waveform_sig_rx =638;
29689: waveform_sig_rx =574;
29690: waveform_sig_rx =942;
29691: waveform_sig_rx =597;
29692: waveform_sig_rx =603;
29693: waveform_sig_rx =1010;
29694: waveform_sig_rx =637;
29695: waveform_sig_rx =603;
29696: waveform_sig_rx =1052;
29697: waveform_sig_rx =619;
29698: waveform_sig_rx =724;
29699: waveform_sig_rx =924;
29700: waveform_sig_rx =784;
29701: waveform_sig_rx =715;
29702: waveform_sig_rx =847;
29703: waveform_sig_rx =902;
29704: waveform_sig_rx =746;
29705: waveform_sig_rx =733;
29706: waveform_sig_rx =991;
29707: waveform_sig_rx =789;
29708: waveform_sig_rx =658;
29709: waveform_sig_rx =1059;
29710: waveform_sig_rx =799;
29711: waveform_sig_rx =688;
29712: waveform_sig_rx =997;
29713: waveform_sig_rx =894;
29714: waveform_sig_rx =723;
29715: waveform_sig_rx =923;
29716: waveform_sig_rx =953;
29717: waveform_sig_rx =799;
29718: waveform_sig_rx =797;
29719: waveform_sig_rx =1056;
29720: waveform_sig_rx =869;
29721: waveform_sig_rx =801;
29722: waveform_sig_rx =1007;
29723: waveform_sig_rx =834;
29724: waveform_sig_rx =968;
29725: waveform_sig_rx =887;
29726: waveform_sig_rx =988;
29727: waveform_sig_rx =746;
29728: waveform_sig_rx =1161;
29729: waveform_sig_rx =827;
29730: waveform_sig_rx =818;
29731: waveform_sig_rx =1178;
29732: waveform_sig_rx =776;
29733: waveform_sig_rx =878;
29734: waveform_sig_rx =1211;
29735: waveform_sig_rx =753;
29736: waveform_sig_rx =881;
29737: waveform_sig_rx =1187;
29738: waveform_sig_rx =806;
29739: waveform_sig_rx =964;
29740: waveform_sig_rx =1038;
29741: waveform_sig_rx =1022;
29742: waveform_sig_rx =841;
29743: waveform_sig_rx =1002;
29744: waveform_sig_rx =1145;
29745: waveform_sig_rx =832;
29746: waveform_sig_rx =954;
29747: waveform_sig_rx =1186;
29748: waveform_sig_rx =877;
29749: waveform_sig_rx =954;
29750: waveform_sig_rx =1181;
29751: waveform_sig_rx =949;
29752: waveform_sig_rx =929;
29753: waveform_sig_rx =1092;
29754: waveform_sig_rx =1108;
29755: waveform_sig_rx =890;
29756: waveform_sig_rx =1041;
29757: waveform_sig_rx =1180;
29758: waveform_sig_rx =914;
29759: waveform_sig_rx =970;
29760: waveform_sig_rx =1261;
29761: waveform_sig_rx =968;
29762: waveform_sig_rx =997;
29763: waveform_sig_rx =1136;
29764: waveform_sig_rx =956;
29765: waveform_sig_rx =1110;
29766: waveform_sig_rx =1048;
29767: waveform_sig_rx =1091;
29768: waveform_sig_rx =910;
29769: waveform_sig_rx =1306;
29770: waveform_sig_rx =902;
29771: waveform_sig_rx =1025;
29772: waveform_sig_rx =1301;
29773: waveform_sig_rx =886;
29774: waveform_sig_rx =1119;
29775: waveform_sig_rx =1247;
29776: waveform_sig_rx =954;
29777: waveform_sig_rx =1030;
29778: waveform_sig_rx =1245;
29779: waveform_sig_rx =1008;
29780: waveform_sig_rx =1001;
29781: waveform_sig_rx =1219;
29782: waveform_sig_rx =1158;
29783: waveform_sig_rx =858;
29784: waveform_sig_rx =1240;
29785: waveform_sig_rx =1192;
29786: waveform_sig_rx =939;
29787: waveform_sig_rx =1124;
29788: waveform_sig_rx =1245;
29789: waveform_sig_rx =1014;
29790: waveform_sig_rx =1035;
29791: waveform_sig_rx =1272;
29792: waveform_sig_rx =1074;
29793: waveform_sig_rx =1011;
29794: waveform_sig_rx =1194;
29795: waveform_sig_rx =1225;
29796: waveform_sig_rx =973;
29797: waveform_sig_rx =1132;
29798: waveform_sig_rx =1307;
29799: waveform_sig_rx =963;
29800: waveform_sig_rx =1073;
29801: waveform_sig_rx =1369;
29802: waveform_sig_rx =983;
29803: waveform_sig_rx =1153;
29804: waveform_sig_rx =1188;
29805: waveform_sig_rx =1021;
29806: waveform_sig_rx =1245;
29807: waveform_sig_rx =1078;
29808: waveform_sig_rx =1187;
29809: waveform_sig_rx =1012;
29810: waveform_sig_rx =1333;
29811: waveform_sig_rx =991;
29812: waveform_sig_rx =1116;
29813: waveform_sig_rx =1294;
29814: waveform_sig_rx =987;
29815: waveform_sig_rx =1122;
29816: waveform_sig_rx =1306;
29817: waveform_sig_rx =1027;
29818: waveform_sig_rx =1035;
29819: waveform_sig_rx =1349;
29820: waveform_sig_rx =1059;
29821: waveform_sig_rx =1029;
29822: waveform_sig_rx =1318;
29823: waveform_sig_rx =1145;
29824: waveform_sig_rx =897;
29825: waveform_sig_rx =1319;
29826: waveform_sig_rx =1153;
29827: waveform_sig_rx =1032;
29828: waveform_sig_rx =1169;
29829: waveform_sig_rx =1250;
29830: waveform_sig_rx =1100;
29831: waveform_sig_rx =1039;
29832: waveform_sig_rx =1305;
29833: waveform_sig_rx =1130;
29834: waveform_sig_rx =1003;
29835: waveform_sig_rx =1254;
29836: waveform_sig_rx =1228;
29837: waveform_sig_rx =956;
29838: waveform_sig_rx =1198;
29839: waveform_sig_rx =1307;
29840: waveform_sig_rx =950;
29841: waveform_sig_rx =1165;
29842: waveform_sig_rx =1345;
29843: waveform_sig_rx =986;
29844: waveform_sig_rx =1221;
29845: waveform_sig_rx =1136;
29846: waveform_sig_rx =1095;
29847: waveform_sig_rx =1243;
29848: waveform_sig_rx =1061;
29849: waveform_sig_rx =1222;
29850: waveform_sig_rx =979;
29851: waveform_sig_rx =1325;
29852: waveform_sig_rx =1017;
29853: waveform_sig_rx =1075;
29854: waveform_sig_rx =1332;
29855: waveform_sig_rx =992;
29856: waveform_sig_rx =1104;
29857: waveform_sig_rx =1345;
29858: waveform_sig_rx =974;
29859: waveform_sig_rx =1035;
29860: waveform_sig_rx =1371;
29861: waveform_sig_rx =973;
29862: waveform_sig_rx =1047;
29863: waveform_sig_rx =1320;
29864: waveform_sig_rx =1046;
29865: waveform_sig_rx =948;
29866: waveform_sig_rx =1269;
29867: waveform_sig_rx =1083;
29868: waveform_sig_rx =1058;
29869: waveform_sig_rx =1086;
29870: waveform_sig_rx =1234;
29871: waveform_sig_rx =1045;
29872: waveform_sig_rx =986;
29873: waveform_sig_rx =1297;
29874: waveform_sig_rx =1048;
29875: waveform_sig_rx =956;
29876: waveform_sig_rx =1238;
29877: waveform_sig_rx =1138;
29878: waveform_sig_rx =909;
29879: waveform_sig_rx =1175;
29880: waveform_sig_rx =1190;
29881: waveform_sig_rx =904;
29882: waveform_sig_rx =1109;
29883: waveform_sig_rx =1227;
29884: waveform_sig_rx =948;
29885: waveform_sig_rx =1138;
29886: waveform_sig_rx =1033;
29887: waveform_sig_rx =1090;
29888: waveform_sig_rx =1124;
29889: waveform_sig_rx =1008;
29890: waveform_sig_rx =1188;
29891: waveform_sig_rx =874;
29892: waveform_sig_rx =1309;
29893: waveform_sig_rx =939;
29894: waveform_sig_rx =987;
29895: waveform_sig_rx =1298;
29896: waveform_sig_rx =846;
29897: waveform_sig_rx =1022;
29898: waveform_sig_rx =1286;
29899: waveform_sig_rx =808;
29900: waveform_sig_rx =1003;
29901: waveform_sig_rx =1248;
29902: waveform_sig_rx =825;
29903: waveform_sig_rx =1005;
29904: waveform_sig_rx =1167;
29905: waveform_sig_rx =973;
29906: waveform_sig_rx =897;
29907: waveform_sig_rx =1139;
29908: waveform_sig_rx =1028;
29909: waveform_sig_rx =916;
29910: waveform_sig_rx =971;
29911: waveform_sig_rx =1191;
29912: waveform_sig_rx =873;
29913: waveform_sig_rx =914;
29914: waveform_sig_rx =1203;
29915: waveform_sig_rx =875;
29916: waveform_sig_rx =876;
29917: waveform_sig_rx =1142;
29918: waveform_sig_rx =978;
29919: waveform_sig_rx =805;
29920: waveform_sig_rx =1074;
29921: waveform_sig_rx =1040;
29922: waveform_sig_rx =823;
29923: waveform_sig_rx =981;
29924: waveform_sig_rx =1075;
29925: waveform_sig_rx =862;
29926: waveform_sig_rx =953;
29927: waveform_sig_rx =914;
29928: waveform_sig_rx =971;
29929: waveform_sig_rx =903;
29930: waveform_sig_rx =942;
29931: waveform_sig_rx =947;
29932: waveform_sig_rx =727;
29933: waveform_sig_rx =1200;
29934: waveform_sig_rx =675;
29935: waveform_sig_rx =898;
29936: waveform_sig_rx =1095;
29937: waveform_sig_rx =626;
29938: waveform_sig_rx =964;
29939: waveform_sig_rx =1051;
29940: waveform_sig_rx =679;
29941: waveform_sig_rx =880;
29942: waveform_sig_rx =1027;
29943: waveform_sig_rx =711;
29944: waveform_sig_rx =821;
29945: waveform_sig_rx =974;
29946: waveform_sig_rx =807;
29947: waveform_sig_rx =693;
29948: waveform_sig_rx =963;
29949: waveform_sig_rx =853;
29950: waveform_sig_rx =742;
29951: waveform_sig_rx =791;
29952: waveform_sig_rx =1014;
29953: waveform_sig_rx =643;
29954: waveform_sig_rx =764;
29955: waveform_sig_rx =1029;
29956: waveform_sig_rx =654;
29957: waveform_sig_rx =745;
29958: waveform_sig_rx =918;
29959: waveform_sig_rx =764;
29960: waveform_sig_rx =690;
29961: waveform_sig_rx =810;
29962: waveform_sig_rx =877;
29963: waveform_sig_rx =619;
29964: waveform_sig_rx =722;
29965: waveform_sig_rx =960;
29966: waveform_sig_rx =591;
29967: waveform_sig_rx =770;
29968: waveform_sig_rx =760;
29969: waveform_sig_rx =706;
29970: waveform_sig_rx =753;
29971: waveform_sig_rx =739;
29972: waveform_sig_rx =684;
29973: waveform_sig_rx =611;
29974: waveform_sig_rx =948;
29975: waveform_sig_rx =460;
29976: waveform_sig_rx =772;
29977: waveform_sig_rx =827;
29978: waveform_sig_rx =467;
29979: waveform_sig_rx =762;
29980: waveform_sig_rx =795;
29981: waveform_sig_rx =484;
29982: waveform_sig_rx =637;
29983: waveform_sig_rx =810;
29984: waveform_sig_rx =491;
29985: waveform_sig_rx =614;
29986: waveform_sig_rx =743;
29987: waveform_sig_rx =604;
29988: waveform_sig_rx =435;
29989: waveform_sig_rx =746;
29990: waveform_sig_rx =629;
29991: waveform_sig_rx =456;
29992: waveform_sig_rx =604;
29993: waveform_sig_rx =737;
29994: waveform_sig_rx =364;
29995: waveform_sig_rx =588;
29996: waveform_sig_rx =702;
29997: waveform_sig_rx =447;
29998: waveform_sig_rx =525;
29999: waveform_sig_rx =607;
30000: waveform_sig_rx =593;
30001: waveform_sig_rx =363;
30002: waveform_sig_rx =596;
30003: waveform_sig_rx =675;
30004: waveform_sig_rx =285;
30005: waveform_sig_rx =560;
30006: waveform_sig_rx =690;
30007: waveform_sig_rx =286;
30008: waveform_sig_rx =604;
30009: waveform_sig_rx =421;
30010: waveform_sig_rx =449;
30011: waveform_sig_rx =517;
30012: waveform_sig_rx =426;
30013: waveform_sig_rx =458;
30014: waveform_sig_rx =359;
30015: waveform_sig_rx =621;
30016: waveform_sig_rx =213;
30017: waveform_sig_rx =476;
30018: waveform_sig_rx =532;
30019: waveform_sig_rx =239;
30020: waveform_sig_rx =495;
30021: waveform_sig_rx =519;
30022: waveform_sig_rx =230;
30023: waveform_sig_rx =379;
30024: waveform_sig_rx =545;
30025: waveform_sig_rx =231;
30026: waveform_sig_rx =297;
30027: waveform_sig_rx =511;
30028: waveform_sig_rx =293;
30029: waveform_sig_rx =159;
30030: waveform_sig_rx =575;
30031: waveform_sig_rx =281;
30032: waveform_sig_rx =222;
30033: waveform_sig_rx =380;
30034: waveform_sig_rx =394;
30035: waveform_sig_rx =208;
30036: waveform_sig_rx =265;
30037: waveform_sig_rx =405;
30038: waveform_sig_rx =222;
30039: waveform_sig_rx =141;
30040: waveform_sig_rx =414;
30041: waveform_sig_rx =290;
30042: waveform_sig_rx =26;
30043: waveform_sig_rx =394;
30044: waveform_sig_rx =293;
30045: waveform_sig_rx =49;
30046: waveform_sig_rx =315;
30047: waveform_sig_rx =326;
30048: waveform_sig_rx =40;
30049: waveform_sig_rx =313;
30050: waveform_sig_rx =121;
30051: waveform_sig_rx =200;
30052: waveform_sig_rx =213;
30053: waveform_sig_rx =129;
30054: waveform_sig_rx =181;
30055: waveform_sig_rx =68;
30056: waveform_sig_rx =307;
30057: waveform_sig_rx =-24;
30058: waveform_sig_rx =160;
30059: waveform_sig_rx =239;
30060: waveform_sig_rx =-61;
30061: waveform_sig_rx =122;
30062: waveform_sig_rx =301;
30063: waveform_sig_rx =-117;
30064: waveform_sig_rx =89;
30065: waveform_sig_rx =319;
30066: waveform_sig_rx =-172;
30067: waveform_sig_rx =91;
30068: waveform_sig_rx =217;
30069: waveform_sig_rx =-70;
30070: waveform_sig_rx =-71;
30071: waveform_sig_rx =219;
30072: waveform_sig_rx =-25;
30073: waveform_sig_rx =-58;
30074: waveform_sig_rx =28;
30075: waveform_sig_rx =128;
30076: waveform_sig_rx =-119;
30077: waveform_sig_rx =-42;
30078: waveform_sig_rx =148;
30079: waveform_sig_rx =-86;
30080: waveform_sig_rx =-152;
30081: waveform_sig_rx =157;
30082: waveform_sig_rx =-55;
30083: waveform_sig_rx =-251;
30084: waveform_sig_rx =128;
30085: waveform_sig_rx =-58;
30086: waveform_sig_rx =-241;
30087: waveform_sig_rx =13;
30088: waveform_sig_rx =4;
30089: waveform_sig_rx =-212;
30090: waveform_sig_rx =-34;
30091: waveform_sig_rx =-190;
30092: waveform_sig_rx =-53;
30093: waveform_sig_rx =-154;
30094: waveform_sig_rx =-120;
30095: waveform_sig_rx =-131;
30096: waveform_sig_rx =-265;
30097: waveform_sig_rx =40;
30098: waveform_sig_rx =-367;
30099: waveform_sig_rx =-165;
30100: waveform_sig_rx =-21;
30101: waveform_sig_rx =-445;
30102: waveform_sig_rx =-134;
30103: waveform_sig_rx =7;
30104: waveform_sig_rx =-490;
30105: waveform_sig_rx =-129;
30106: waveform_sig_rx =-49;
30107: waveform_sig_rx =-490;
30108: waveform_sig_rx =-165;
30109: waveform_sig_rx =-156;
30110: waveform_sig_rx =-336;
30111: waveform_sig_rx =-359;
30112: waveform_sig_rx =-125;
30113: waveform_sig_rx =-304;
30114: waveform_sig_rx =-377;
30115: waveform_sig_rx =-280;
30116: waveform_sig_rx =-171;
30117: waveform_sig_rx =-454;
30118: waveform_sig_rx =-320;
30119: waveform_sig_rx =-141;
30120: waveform_sig_rx =-450;
30121: waveform_sig_rx =-422;
30122: waveform_sig_rx =-116;
30123: waveform_sig_rx =-418;
30124: waveform_sig_rx =-483;
30125: waveform_sig_rx =-168;
30126: waveform_sig_rx =-403;
30127: waveform_sig_rx =-452;
30128: waveform_sig_rx =-361;
30129: waveform_sig_rx =-282;
30130: waveform_sig_rx =-503;
30131: waveform_sig_rx =-401;
30132: waveform_sig_rx =-406;
30133: waveform_sig_rx =-389;
30134: waveform_sig_rx =-478;
30135: waveform_sig_rx =-350;
30136: waveform_sig_rx =-514;
30137: waveform_sig_rx =-515;
30138: waveform_sig_rx =-228;
30139: waveform_sig_rx =-712;
30140: waveform_sig_rx =-379;
30141: waveform_sig_rx =-351;
30142: waveform_sig_rx =-725;
30143: waveform_sig_rx =-372;
30144: waveform_sig_rx =-366;
30145: waveform_sig_rx =-783;
30146: waveform_sig_rx =-417;
30147: waveform_sig_rx =-396;
30148: waveform_sig_rx =-743;
30149: waveform_sig_rx =-445;
30150: waveform_sig_rx =-483;
30151: waveform_sig_rx =-603;
30152: waveform_sig_rx =-668;
30153: waveform_sig_rx =-435;
30154: waveform_sig_rx =-545;
30155: waveform_sig_rx =-710;
30156: waveform_sig_rx =-543;
30157: waveform_sig_rx =-430;
30158: waveform_sig_rx =-819;
30159: waveform_sig_rx =-553;
30160: waveform_sig_rx =-460;
30161: waveform_sig_rx =-783;
30162: waveform_sig_rx =-635;
30163: waveform_sig_rx =-486;
30164: waveform_sig_rx =-689;
30165: waveform_sig_rx =-758;
30166: waveform_sig_rx =-557;
30167: waveform_sig_rx =-615;
30168: waveform_sig_rx =-795;
30169: waveform_sig_rx =-647;
30170: waveform_sig_rx =-505;
30171: waveform_sig_rx =-864;
30172: waveform_sig_rx =-612;
30173: waveform_sig_rx =-725;
30174: waveform_sig_rx =-695;
30175: waveform_sig_rx =-712;
30176: waveform_sig_rx =-640;
30177: waveform_sig_rx =-806;
30178: waveform_sig_rx =-737;
30179: waveform_sig_rx =-564;
30180: waveform_sig_rx =-1002;
30181: waveform_sig_rx =-618;
30182: waveform_sig_rx =-668;
30183: waveform_sig_rx =-992;
30184: waveform_sig_rx =-594;
30185: waveform_sig_rx =-665;
30186: waveform_sig_rx =-1002;
30187: waveform_sig_rx =-636;
30188: waveform_sig_rx =-709;
30189: waveform_sig_rx =-946;
30190: waveform_sig_rx =-740;
30191: waveform_sig_rx =-715;
30192: waveform_sig_rx =-808;
30193: waveform_sig_rx =-984;
30194: waveform_sig_rx =-616;
30195: waveform_sig_rx =-845;
30196: waveform_sig_rx =-1000;
30197: waveform_sig_rx =-713;
30198: waveform_sig_rx =-756;
30199: waveform_sig_rx =-1033;
30200: waveform_sig_rx =-748;
30201: waveform_sig_rx =-761;
30202: waveform_sig_rx =-949;
30203: waveform_sig_rx =-907;
30204: waveform_sig_rx =-727;
30205: waveform_sig_rx =-881;
30206: waveform_sig_rx =-1012;
30207: waveform_sig_rx =-712;
30208: waveform_sig_rx =-817;
30209: waveform_sig_rx =-1045;
30210: waveform_sig_rx =-809;
30211: waveform_sig_rx =-751;
30212: waveform_sig_rx =-1080;
30213: waveform_sig_rx =-791;
30214: waveform_sig_rx =-953;
30215: waveform_sig_rx =-880;
30216: waveform_sig_rx =-898;
30217: waveform_sig_rx =-881;
30218: waveform_sig_rx =-1031;
30219: waveform_sig_rx =-904;
30220: waveform_sig_rx =-814;
30221: waveform_sig_rx =-1169;
30222: waveform_sig_rx =-786;
30223: waveform_sig_rx =-938;
30224: waveform_sig_rx =-1141;
30225: waveform_sig_rx =-841;
30226: waveform_sig_rx =-895;
30227: waveform_sig_rx =-1147;
30228: waveform_sig_rx =-904;
30229: waveform_sig_rx =-853;
30230: waveform_sig_rx =-1134;
30231: waveform_sig_rx =-988;
30232: waveform_sig_rx =-846;
30233: waveform_sig_rx =-1097;
30234: waveform_sig_rx =-1143;
30235: waveform_sig_rx =-764;
30236: waveform_sig_rx =-1123;
30237: waveform_sig_rx =-1114;
30238: waveform_sig_rx =-923;
30239: waveform_sig_rx =-975;
30240: waveform_sig_rx =-1161;
30241: waveform_sig_rx =-986;
30242: waveform_sig_rx =-923;
30243: waveform_sig_rx =-1127;
30244: waveform_sig_rx =-1103;
30245: waveform_sig_rx =-880;
30246: waveform_sig_rx =-1093;
30247: waveform_sig_rx =-1208;
30248: waveform_sig_rx =-896;
30249: waveform_sig_rx =-1057;
30250: waveform_sig_rx =-1248;
30251: waveform_sig_rx =-966;
30252: waveform_sig_rx =-975;
30253: waveform_sig_rx =-1273;
30254: waveform_sig_rx =-948;
30255: waveform_sig_rx =-1189;
30256: waveform_sig_rx =-1045;
30257: waveform_sig_rx =-1083;
30258: waveform_sig_rx =-1080;
30259: waveform_sig_rx =-1155;
30260: waveform_sig_rx =-1078;
30261: waveform_sig_rx =-1005;
30262: waveform_sig_rx =-1271;
30263: waveform_sig_rx =-991;
30264: waveform_sig_rx =-1060;
30265: waveform_sig_rx =-1266;
30266: waveform_sig_rx =-1015;
30267: waveform_sig_rx =-978;
30268: waveform_sig_rx =-1349;
30269: waveform_sig_rx =-1005;
30270: waveform_sig_rx =-971;
30271: waveform_sig_rx =-1346;
30272: waveform_sig_rx =-1028;
30273: waveform_sig_rx =-1004;
30274: waveform_sig_rx =-1273;
30275: waveform_sig_rx =-1188;
30276: waveform_sig_rx =-940;
30277: waveform_sig_rx =-1243;
30278: waveform_sig_rx =-1194;
30279: waveform_sig_rx =-1080;
30280: waveform_sig_rx =-1066;
30281: waveform_sig_rx =-1277;
30282: waveform_sig_rx =-1123;
30283: waveform_sig_rx =-1034;
30284: waveform_sig_rx =-1253;
30285: waveform_sig_rx =-1223;
30286: waveform_sig_rx =-935;
30287: waveform_sig_rx =-1226;
30288: waveform_sig_rx =-1293;
30289: waveform_sig_rx =-918;
30290: waveform_sig_rx =-1214;
30291: waveform_sig_rx =-1285;
30292: waveform_sig_rx =-1006;
30293: waveform_sig_rx =-1106;
30294: waveform_sig_rx =-1274;
30295: waveform_sig_rx =-1022;
30296: waveform_sig_rx =-1261;
30297: waveform_sig_rx =-1042;
30298: waveform_sig_rx =-1236;
30299: waveform_sig_rx =-1103;
30300: waveform_sig_rx =-1214;
30301: waveform_sig_rx =-1177;
30302: waveform_sig_rx =-1014;
30303: waveform_sig_rx =-1370;
30304: waveform_sig_rx =-1034;
30305: waveform_sig_rx =-1074;
30306: waveform_sig_rx =-1384;
30307: waveform_sig_rx =-1019;
30308: waveform_sig_rx =-1048;
30309: waveform_sig_rx =-1430;
30310: waveform_sig_rx =-1001;
30311: waveform_sig_rx =-1066;
30312: waveform_sig_rx =-1396;
30313: waveform_sig_rx =-1033;
30314: waveform_sig_rx =-1054;
30315: waveform_sig_rx =-1313;
30316: waveform_sig_rx =-1191;
30317: waveform_sig_rx =-1036;
30318: waveform_sig_rx =-1251;
30319: waveform_sig_rx =-1209;
30320: waveform_sig_rx =-1140;
30321: waveform_sig_rx =-1045;
30322: waveform_sig_rx =-1350;
30323: waveform_sig_rx =-1107;
30324: waveform_sig_rx =-1008;
30325: waveform_sig_rx =-1349;
30326: waveform_sig_rx =-1182;
30327: waveform_sig_rx =-979;
30328: waveform_sig_rx =-1300;
30329: waveform_sig_rx =-1256;
30330: waveform_sig_rx =-983;
30331: waveform_sig_rx =-1217;
30332: waveform_sig_rx =-1268;
30333: waveform_sig_rx =-1046;
30334: waveform_sig_rx =-1122;
30335: waveform_sig_rx =-1265;
30336: waveform_sig_rx =-1086;
30337: waveform_sig_rx =-1251;
30338: waveform_sig_rx =-1037;
30339: waveform_sig_rx =-1262;
30340: waveform_sig_rx =-1026;
30341: waveform_sig_rx =-1259;
30342: waveform_sig_rx =-1148;
30343: waveform_sig_rx =-979;
30344: waveform_sig_rx =-1419;
30345: waveform_sig_rx =-972;
30346: waveform_sig_rx =-1068;
30347: waveform_sig_rx =-1397;
30348: waveform_sig_rx =-893;
30349: waveform_sig_rx =-1099;
30350: waveform_sig_rx =-1376;
30351: waveform_sig_rx =-932;
30352: waveform_sig_rx =-1096;
30353: waveform_sig_rx =-1299;
30354: waveform_sig_rx =-999;
30355: waveform_sig_rx =-1072;
30356: waveform_sig_rx =-1252;
30357: waveform_sig_rx =-1154;
30358: waveform_sig_rx =-980;
30359: waveform_sig_rx =-1163;
30360: waveform_sig_rx =-1200;
30361: waveform_sig_rx =-1045;
30362: waveform_sig_rx =-995;
30363: waveform_sig_rx =-1336;
30364: waveform_sig_rx =-982;
30365: waveform_sig_rx =-982;
30366: waveform_sig_rx =-1303;
30367: waveform_sig_rx =-1042;
30368: waveform_sig_rx =-951;
30369: waveform_sig_rx =-1219;
30370: waveform_sig_rx =-1120;
30371: waveform_sig_rx =-959;
30372: waveform_sig_rx =-1120;
30373: waveform_sig_rx =-1177;
30374: waveform_sig_rx =-988;
30375: waveform_sig_rx =-986;
30376: waveform_sig_rx =-1209;
30377: waveform_sig_rx =-1008;
30378: waveform_sig_rx =-1141;
30379: waveform_sig_rx =-991;
30380: waveform_sig_rx =-1156;
30381: waveform_sig_rx =-899;
30382: waveform_sig_rx =-1241;
30383: waveform_sig_rx =-975;
30384: waveform_sig_rx =-920;
30385: waveform_sig_rx =-1338;
30386: waveform_sig_rx =-763;
30387: waveform_sig_rx =-1081;
30388: waveform_sig_rx =-1225;
30389: waveform_sig_rx =-778;
30390: waveform_sig_rx =-1096;
30391: waveform_sig_rx =-1175;
30392: waveform_sig_rx =-868;
30393: waveform_sig_rx =-994;
30394: waveform_sig_rx =-1139;
30395: waveform_sig_rx =-954;
30396: waveform_sig_rx =-905;
30397: waveform_sig_rx =-1127;
30398: waveform_sig_rx =-1017;
30399: waveform_sig_rx =-828;
30400: waveform_sig_rx =-1062;
30401: waveform_sig_rx =-1067;
30402: waveform_sig_rx =-872;
30403: waveform_sig_rx =-859;
30404: waveform_sig_rx =-1211;
30405: waveform_sig_rx =-804;
30406: waveform_sig_rx =-887;
30407: waveform_sig_rx =-1154;
30408: waveform_sig_rx =-846;
30409: waveform_sig_rx =-875;
30410: waveform_sig_rx =-1005;
30411: waveform_sig_rx =-984;
30412: waveform_sig_rx =-835;
30413: waveform_sig_rx =-871;
30414: waveform_sig_rx =-1110;
30415: waveform_sig_rx =-794;
30416: waveform_sig_rx =-825;
30417: waveform_sig_rx =-1130;
30418: waveform_sig_rx =-739;
30419: waveform_sig_rx =-995;
30420: waveform_sig_rx =-843;
30421: waveform_sig_rx =-906;
30422: waveform_sig_rx =-812;
30423: waveform_sig_rx =-1042;
30424: waveform_sig_rx =-732;
30425: waveform_sig_rx =-840;
30426: waveform_sig_rx =-1079;
30427: waveform_sig_rx =-631;
30428: waveform_sig_rx =-951;
30429: waveform_sig_rx =-1000;
30430: waveform_sig_rx =-658;
30431: waveform_sig_rx =-891;
30432: waveform_sig_rx =-978;
30433: waveform_sig_rx =-697;
30434: waveform_sig_rx =-799;
30435: waveform_sig_rx =-948;
30436: waveform_sig_rx =-758;
30437: waveform_sig_rx =-690;
30438: waveform_sig_rx =-938;
30439: waveform_sig_rx =-845;
30440: waveform_sig_rx =-603;
30441: waveform_sig_rx =-906;
30442: waveform_sig_rx =-869;
30443: waveform_sig_rx =-617;
30444: waveform_sig_rx =-772;
30445: waveform_sig_rx =-939;
30446: waveform_sig_rx =-605;
30447: waveform_sig_rx =-762;
30448: waveform_sig_rx =-831;
30449: waveform_sig_rx =-723;
30450: waveform_sig_rx =-620;
30451: waveform_sig_rx =-761;
30452: waveform_sig_rx =-874;
30453: waveform_sig_rx =-512;
30454: waveform_sig_rx =-761;
30455: waveform_sig_rx =-895;
30456: waveform_sig_rx =-471;
30457: waveform_sig_rx =-698;
30458: waveform_sig_rx =-819;
30459: waveform_sig_rx =-535;
30460: waveform_sig_rx =-842;
30461: waveform_sig_rx =-540;
30462: waveform_sig_rx =-723;
30463: waveform_sig_rx =-595;
30464: waveform_sig_rx =-784;
30465: waveform_sig_rx =-551;
30466: waveform_sig_rx =-622;
30467: waveform_sig_rx =-826;
30468: waveform_sig_rx =-446;
30469: waveform_sig_rx =-692;
30470: waveform_sig_rx =-749;
30471: waveform_sig_rx =-435;
30472: waveform_sig_rx =-647;
30473: waveform_sig_rx =-750;
30474: waveform_sig_rx =-461;
30475: waveform_sig_rx =-544;
30476: waveform_sig_rx =-750;
30477: waveform_sig_rx =-524;
30478: waveform_sig_rx =-412;
30479: waveform_sig_rx =-783;
30480: waveform_sig_rx =-545;
30481: waveform_sig_rx =-367;
30482: waveform_sig_rx =-731;
30483: waveform_sig_rx =-554;
30484: waveform_sig_rx =-450;
30485: waveform_sig_rx =-524;
30486: waveform_sig_rx =-625;
30487: waveform_sig_rx =-437;
30488: waveform_sig_rx =-432;
30489: waveform_sig_rx =-616;
30490: waveform_sig_rx =-518;
30491: waveform_sig_rx =-294;
30492: waveform_sig_rx =-617;
30493: waveform_sig_rx =-559;
30494: waveform_sig_rx =-238;
30495: waveform_sig_rx =-575;
30496: waveform_sig_rx =-555;
30497: waveform_sig_rx =-260;
30498: waveform_sig_rx =-468;
30499: waveform_sig_rx =-533;
30500: waveform_sig_rx =-328;
30501: waveform_sig_rx =-549;
30502: waveform_sig_rx =-289;
30503: waveform_sig_rx =-492;
30504: waveform_sig_rx =-304;
30505: waveform_sig_rx =-532;
30506: waveform_sig_rx =-292;
30507: waveform_sig_rx =-357;
30508: waveform_sig_rx =-546;
30509: waveform_sig_rx =-196;
30510: waveform_sig_rx =-419;
30511: waveform_sig_rx =-491;
30512: waveform_sig_rx =-185;
30513: waveform_sig_rx =-307;
30514: waveform_sig_rx =-556;
30515: waveform_sig_rx =-149;
30516: waveform_sig_rx =-265;
30517: waveform_sig_rx =-547;
30518: waveform_sig_rx =-135;
30519: waveform_sig_rx =-230;
30520: waveform_sig_rx =-507;
30521: waveform_sig_rx =-187;
30522: waveform_sig_rx =-205;
30523: waveform_sig_rx =-370;
30524: waveform_sig_rx =-297;
30525: waveform_sig_rx =-211;
30526: waveform_sig_rx =-162;
30527: waveform_sig_rx =-442;
30528: waveform_sig_rx =-116;
30529: waveform_sig_rx =-139;
30530: waveform_sig_rx =-402;
30531: waveform_sig_rx =-168;
30532: waveform_sig_rx =-57;
30533: waveform_sig_rx =-357;
30534: waveform_sig_rx =-225;
30535: waveform_sig_rx =14;
30536: waveform_sig_rx =-296;
30537: waveform_sig_rx =-254;
30538: waveform_sig_rx =15;
30539: waveform_sig_rx =-202;
30540: waveform_sig_rx =-189;
30541: waveform_sig_rx =-76;
30542: waveform_sig_rx =-234;
30543: waveform_sig_rx =19;
30544: waveform_sig_rx =-237;
30545: waveform_sig_rx =23;
30546: waveform_sig_rx =-265;
30547: waveform_sig_rx =-7;
30548: waveform_sig_rx =-28;
30549: waveform_sig_rx =-298;
30550: waveform_sig_rx =130;
30551: waveform_sig_rx =-103;
30552: waveform_sig_rx =-262;
30553: waveform_sig_rx =194;
30554: waveform_sig_rx =-101;
30555: waveform_sig_rx =-250;
30556: waveform_sig_rx =206;
30557: waveform_sig_rx =-81;
30558: waveform_sig_rx =-169;
30559: waveform_sig_rx =144;
30560: waveform_sig_rx =13;
30561: waveform_sig_rx =-141;
30562: waveform_sig_rx =53;
30563: waveform_sig_rx =109;
30564: waveform_sig_rx =-45;
30565: waveform_sig_rx =-55;
30566: waveform_sig_rx =146;
30567: waveform_sig_rx =104;
30568: waveform_sig_rx =-156;
30569: waveform_sig_rx =227;
30570: waveform_sig_rx =98;
30571: waveform_sig_rx =-122;
30572: waveform_sig_rx =138;
30573: waveform_sig_rx =195;
30574: waveform_sig_rx =-63;
30575: waveform_sig_rx =94;
30576: waveform_sig_rx =240;
30577: waveform_sig_rx =29;
30578: waveform_sig_rx =63;
30579: waveform_sig_rx =248;
30580: waveform_sig_rx =144;
30581: waveform_sig_rx =56;
30582: waveform_sig_rx =202;
30583: waveform_sig_rx =108;
30584: waveform_sig_rx =222;
30585: waveform_sig_rx =90;
30586: waveform_sig_rx =338;
30587: waveform_sig_rx =-33;
30588: waveform_sig_rx =374;
30589: waveform_sig_rx =202;
30590: waveform_sig_rx =-1;
30591: waveform_sig_rx =486;
30592: waveform_sig_rx =114;
30593: waveform_sig_rx =88;
30594: waveform_sig_rx =497;
30595: waveform_sig_rx =127;
30596: waveform_sig_rx =114;
30597: waveform_sig_rx =469;
30598: waveform_sig_rx =191;
30599: waveform_sig_rx =167;
30600: waveform_sig_rx =386;
30601: waveform_sig_rx =326;
30602: waveform_sig_rx =165;
30603: waveform_sig_rx =317;
30604: waveform_sig_rx =453;
30605: waveform_sig_rx =216;
30606: waveform_sig_rx =227;
30607: waveform_sig_rx =494;
30608: waveform_sig_rx =324;
30609: waveform_sig_rx =154;
30610: waveform_sig_rx =550;
30611: waveform_sig_rx =342;
30612: waveform_sig_rx =218;
30613: waveform_sig_rx =476;
30614: waveform_sig_rx =464;
30615: waveform_sig_rx =254;
30616: waveform_sig_rx =381;
30617: waveform_sig_rx =525;
30618: waveform_sig_rx =348;
30619: waveform_sig_rx =283;
30620: waveform_sig_rx =567;
30621: waveform_sig_rx =436;
30622: waveform_sig_rx =274;
30623: waveform_sig_rx =560;
30624: waveform_sig_rx =362;
30625: waveform_sig_rx =493;
30626: waveform_sig_rx =447;
30627: waveform_sig_rx =529;
30628: waveform_sig_rx =287;
30629: waveform_sig_rx =688;
30630: waveform_sig_rx =392;
30631: waveform_sig_rx =364;
30632: waveform_sig_rx =735;
30633: waveform_sig_rx =357;
30634: waveform_sig_rx =421;
30635: waveform_sig_rx =723;
30636: waveform_sig_rx =427;
30637: waveform_sig_rx =385;
30638: waveform_sig_rx =742;
30639: waveform_sig_rx =467;
30640: waveform_sig_rx =459;
30641: waveform_sig_rx =624;
30642: waveform_sig_rx =639;
30643: waveform_sig_rx =413;
30644: waveform_sig_rx =562;
30645: waveform_sig_rx =776;
30646: waveform_sig_rx =422;
30647: waveform_sig_rx =555;
30648: waveform_sig_rx =781;
30649: waveform_sig_rx =504;
30650: waveform_sig_rx =518;
30651: waveform_sig_rx =764;
30652: waveform_sig_rx =604;
30653: waveform_sig_rx =526;
30654: waveform_sig_rx =657;
30655: waveform_sig_rx =787;
30656: waveform_sig_rx =490;
30657: waveform_sig_rx =605;
30658: waveform_sig_rx =832;
30659: waveform_sig_rx =544;
30660: waveform_sig_rx =561;
30661: waveform_sig_rx =844;
30662: waveform_sig_rx =630;
30663: waveform_sig_rx =559;
30664: waveform_sig_rx =794;
30665: waveform_sig_rx =582;
30666: waveform_sig_rx =763;
30667: waveform_sig_rx =696;
30668: waveform_sig_rx =739;
30669: waveform_sig_rx =571;
30670: waveform_sig_rx =913;
30671: waveform_sig_rx =608;
30672: waveform_sig_rx =676;
30673: waveform_sig_rx =904;
30674: waveform_sig_rx =624;
30675: waveform_sig_rx =708;
30676: waveform_sig_rx =915;
30677: waveform_sig_rx =726;
30678: waveform_sig_rx =605;
30679: waveform_sig_rx =999;
30680: waveform_sig_rx =738;
30681: waveform_sig_rx =651;
30682: waveform_sig_rx =915;
30683: waveform_sig_rx =862;
30684: waveform_sig_rx =592;
30685: waveform_sig_rx =880;
30686: waveform_sig_rx =953;
30687: waveform_sig_rx =634;
30688: waveform_sig_rx =817;
30689: waveform_sig_rx =962;
30690: waveform_sig_rx =752;
30691: waveform_sig_rx =773;
30692: waveform_sig_rx =944;
30693: waveform_sig_rx =865;
30694: waveform_sig_rx =726;
30695: waveform_sig_rx =876;
30696: waveform_sig_rx =1031;
30697: waveform_sig_rx =669;
30698: waveform_sig_rx =863;
30699: waveform_sig_rx =1068;
30700: waveform_sig_rx =733;
30701: waveform_sig_rx =833;
30702: waveform_sig_rx =1076;
30703: waveform_sig_rx =814;
30704: waveform_sig_rx =846;
30705: waveform_sig_rx =984;
30706: waveform_sig_rx =790;
30707: waveform_sig_rx =1040;
30708: waveform_sig_rx =858;
30709: waveform_sig_rx =968;
30710: waveform_sig_rx =799;
30711: waveform_sig_rx =1059;
30712: waveform_sig_rx =855;
30713: waveform_sig_rx =853;
30714: waveform_sig_rx =1104;
30715: waveform_sig_rx =872;
30716: waveform_sig_rx =839;
30717: waveform_sig_rx =1156;
30718: waveform_sig_rx =899;
30719: waveform_sig_rx =775;
30720: waveform_sig_rx =1234;
30721: waveform_sig_rx =859;
30722: waveform_sig_rx =844;
30723: waveform_sig_rx =1164;
30724: waveform_sig_rx =981;
30725: waveform_sig_rx =779;
30726: waveform_sig_rx =1072;
30727: waveform_sig_rx =1053;
30728: waveform_sig_rx =857;
30729: waveform_sig_rx =976;
30730: waveform_sig_rx =1077;
30731: waveform_sig_rx =950;
30732: waveform_sig_rx =909;
30733: waveform_sig_rx =1118;
30734: waveform_sig_rx =1047;
30735: waveform_sig_rx =854;
30736: waveform_sig_rx =1086;
30737: waveform_sig_rx =1171;
30738: waveform_sig_rx =777;
30739: waveform_sig_rx =1080;
30740: waveform_sig_rx =1178;
30741: waveform_sig_rx =849;
30742: waveform_sig_rx =1033;
30743: waveform_sig_rx =1176;
30744: waveform_sig_rx =952;
30745: waveform_sig_rx =1047;
30746: waveform_sig_rx =1056;
30747: waveform_sig_rx =994;
30748: waveform_sig_rx =1148;
30749: waveform_sig_rx =948;
30750: waveform_sig_rx =1190;
30751: waveform_sig_rx =891;
30752: waveform_sig_rx =1229;
30753: waveform_sig_rx =1029;
30754: waveform_sig_rx =927;
30755: waveform_sig_rx =1279;
30756: waveform_sig_rx =967;
30757: waveform_sig_rx =961;
30758: waveform_sig_rx =1340;
30759: waveform_sig_rx =968;
30760: waveform_sig_rx =941;
30761: waveform_sig_rx =1373;
30762: waveform_sig_rx =961;
30763: waveform_sig_rx =1011;
30764: waveform_sig_rx =1294;
30765: waveform_sig_rx =1083;
30766: waveform_sig_rx =947;
30767: waveform_sig_rx =1226;
30768: waveform_sig_rx =1154;
30769: waveform_sig_rx =1030;
30770: waveform_sig_rx =1077;
30771: waveform_sig_rx =1227;
30772: waveform_sig_rx =1094;
30773: waveform_sig_rx =961;
30774: waveform_sig_rx =1311;
30775: waveform_sig_rx =1112;
30776: waveform_sig_rx =919;
30777: waveform_sig_rx =1267;
30778: waveform_sig_rx =1181;
30779: waveform_sig_rx =919;
30780: waveform_sig_rx =1230;
30781: waveform_sig_rx =1218;
30782: waveform_sig_rx =1013;
30783: waveform_sig_rx =1113;
30784: waveform_sig_rx =1273;
30785: waveform_sig_rx =1086;
30786: waveform_sig_rx =1091;
30787: waveform_sig_rx =1166;
30788: waveform_sig_rx =1106;
30789: waveform_sig_rx =1176;
30790: waveform_sig_rx =1074;
30791: waveform_sig_rx =1212;
30792: waveform_sig_rx =941;
30793: waveform_sig_rx =1353;
30794: waveform_sig_rx =1019;
30795: waveform_sig_rx =1012;
30796: waveform_sig_rx =1392;
30797: waveform_sig_rx =965;
30798: waveform_sig_rx =1079;
30799: waveform_sig_rx =1414;
30800: waveform_sig_rx =935;
30801: waveform_sig_rx =1083;
30802: waveform_sig_rx =1389;
30803: waveform_sig_rx =964;
30804: waveform_sig_rx =1127;
30805: waveform_sig_rx =1258;
30806: waveform_sig_rx =1138;
30807: waveform_sig_rx =1005;
30808: waveform_sig_rx =1206;
30809: waveform_sig_rx =1231;
30810: waveform_sig_rx =1035;
30811: waveform_sig_rx =1092;
30812: waveform_sig_rx =1316;
30813: waveform_sig_rx =1056;
30814: waveform_sig_rx =1020;
30815: waveform_sig_rx =1361;
30816: waveform_sig_rx =1090;
30817: waveform_sig_rx =1022;
30818: waveform_sig_rx =1297;
30819: waveform_sig_rx =1168;
30820: waveform_sig_rx =988;
30821: waveform_sig_rx =1216;
30822: waveform_sig_rx =1234;
30823: waveform_sig_rx =1038;
30824: waveform_sig_rx =1078;
30825: waveform_sig_rx =1294;
30826: waveform_sig_rx =1080;
30827: waveform_sig_rx =1076;
30828: waveform_sig_rx =1194;
30829: waveform_sig_rx =1082;
30830: waveform_sig_rx =1169;
30831: waveform_sig_rx =1115;
30832: waveform_sig_rx =1185;
30833: waveform_sig_rx =939;
30834: waveform_sig_rx =1389;
30835: waveform_sig_rx =938;
30836: waveform_sig_rx =1073;
30837: waveform_sig_rx =1361;
30838: waveform_sig_rx =881;
30839: waveform_sig_rx =1147;
30840: waveform_sig_rx =1319;
30841: waveform_sig_rx =939;
30842: waveform_sig_rx =1106;
30843: waveform_sig_rx =1289;
30844: waveform_sig_rx =1008;
30845: waveform_sig_rx =1070;
30846: waveform_sig_rx =1224;
30847: waveform_sig_rx =1169;
30848: waveform_sig_rx =929;
30849: waveform_sig_rx =1236;
30850: waveform_sig_rx =1199;
30851: waveform_sig_rx =970;
30852: waveform_sig_rx =1119;
30853: waveform_sig_rx =1268;
30854: waveform_sig_rx =1007;
30855: waveform_sig_rx =1031;
30856: waveform_sig_rx =1295;
30857: waveform_sig_rx =1034;
30858: waveform_sig_rx =1006;
30859: waveform_sig_rx =1210;
30860: waveform_sig_rx =1107;
30861: waveform_sig_rx =960;
30862: waveform_sig_rx =1107;
30863: waveform_sig_rx =1200;
30864: waveform_sig_rx =980;
30865: waveform_sig_rx =985;
30866: waveform_sig_rx =1309;
30867: waveform_sig_rx =950;
30868: waveform_sig_rx =1030;
30869: waveform_sig_rx =1133;
30870: waveform_sig_rx =955;
30871: waveform_sig_rx =1145;
30872: waveform_sig_rx =1053;
30873: waveform_sig_rx =1050;
30874: waveform_sig_rx =950;
30875: waveform_sig_rx =1270;
30876: waveform_sig_rx =838;
30877: waveform_sig_rx =1076;
30878: waveform_sig_rx =1192;
30879: waveform_sig_rx =856;
30880: waveform_sig_rx =1075;
30881: waveform_sig_rx =1188;
30882: waveform_sig_rx =903;
30883: waveform_sig_rx =976;
30884: waveform_sig_rx =1219;
30885: waveform_sig_rx =904;
30886: waveform_sig_rx =945;
30887: waveform_sig_rx =1154;
30888: waveform_sig_rx =1025;
30889: waveform_sig_rx =818;
30890: waveform_sig_rx =1159;
30891: waveform_sig_rx =1047;
30892: waveform_sig_rx =870;
30893: waveform_sig_rx =1032;
30894: waveform_sig_rx =1137;
30895: waveform_sig_rx =845;
30896: waveform_sig_rx =963;
30897: waveform_sig_rx =1124;
30898: waveform_sig_rx =898;
30899: waveform_sig_rx =911;
30900: waveform_sig_rx =1030;
30901: waveform_sig_rx =1075;
30902: waveform_sig_rx =805;
30903: waveform_sig_rx =978;
30904: waveform_sig_rx =1170;
30905: waveform_sig_rx =737;
30906: waveform_sig_rx =966;
30907: waveform_sig_rx =1172;
30908: waveform_sig_rx =731;
30909: waveform_sig_rx =1046;
30910: waveform_sig_rx =903;
30911: waveform_sig_rx =863;
30912: waveform_sig_rx =1036;
30913: waveform_sig_rx =845;
30914: waveform_sig_rx =971;
30915: waveform_sig_rx =789;
30916: waveform_sig_rx =1106;
30917: waveform_sig_rx =749;
30918: waveform_sig_rx =892;
30919: waveform_sig_rx =1066;
30920: waveform_sig_rx =699;
30921: waveform_sig_rx =905;
30922: waveform_sig_rx =1044;
30923: waveform_sig_rx =723;
30924: waveform_sig_rx =827;
30925: waveform_sig_rx =1058;
30926: waveform_sig_rx =774;
30927: waveform_sig_rx =762;
30928: waveform_sig_rx =1028;
30929: waveform_sig_rx =846;
30930: waveform_sig_rx =619;
30931: waveform_sig_rx =1077;
30932: waveform_sig_rx =801;
30933: waveform_sig_rx =729;
30934: waveform_sig_rx =877;
30935: waveform_sig_rx =910;
30936: waveform_sig_rx =766;
30937: waveform_sig_rx =742;
30938: waveform_sig_rx =951;
30939: waveform_sig_rx =784;
30940: waveform_sig_rx =653;
30941: waveform_sig_rx =934;
30942: waveform_sig_rx =866;
30943: waveform_sig_rx =562;
30944: waveform_sig_rx =892;
30945: waveform_sig_rx =893;
30946: waveform_sig_rx =556;
30947: waveform_sig_rx =811;
30948: waveform_sig_rx =884;
30949: waveform_sig_rx =588;
30950: waveform_sig_rx =820;
30951: waveform_sig_rx =681;
30952: waveform_sig_rx =732;
30953: waveform_sig_rx =776;
30954: waveform_sig_rx =662;
30955: waveform_sig_rx =786;
30956: waveform_sig_rx =561;
30957: waveform_sig_rx =930;
30958: waveform_sig_rx =520;
30959: waveform_sig_rx =682;
30960: waveform_sig_rx =839;
30961: waveform_sig_rx =496;
30962: waveform_sig_rx =694;
30963: waveform_sig_rx =854;
30964: waveform_sig_rx =516;
30965: waveform_sig_rx =580;
30966: waveform_sig_rx =890;
30967: waveform_sig_rx =489;
30968: waveform_sig_rx =556;
30969: waveform_sig_rx =853;
30970: waveform_sig_rx =523;
30971: waveform_sig_rx =499;
30972: waveform_sig_rx =825;
30973: waveform_sig_rx =521;
30974: waveform_sig_rx =589;
30975: waveform_sig_rx =554;
30976: waveform_sig_rx =720;
30977: waveform_sig_rx =527;
30978: waveform_sig_rx =438;
30979: waveform_sig_rx =813;
30980: waveform_sig_rx =471;
30981: waveform_sig_rx =429;
30982: waveform_sig_rx =745;
30983: waveform_sig_rx =529;
30984: waveform_sig_rx =384;
30985: waveform_sig_rx =648;
30986: waveform_sig_rx =588;
30987: waveform_sig_rx =357;
30988: waveform_sig_rx =535;
30989: waveform_sig_rx =646;
30990: waveform_sig_rx =345;
30991: waveform_sig_rx =570;
30992: waveform_sig_rx =406;
30993: waveform_sig_rx =503;
30994: waveform_sig_rx =482;
30995: waveform_sig_rx =411;
30996: waveform_sig_rx =531;
30997: waveform_sig_rx =271;
30998: waveform_sig_rx =674;
30999: waveform_sig_rx =285;
31000: waveform_sig_rx =394;
31001: waveform_sig_rx =647;
31002: waveform_sig_rx =182;
31003: waveform_sig_rx =412;
31004: waveform_sig_rx =632;
31005: waveform_sig_rx =114;
31006: waveform_sig_rx =414;
31007: waveform_sig_rx =581;
31008: waveform_sig_rx =140;
31009: waveform_sig_rx =408;
31010: waveform_sig_rx =467;
31011: waveform_sig_rx =288;
31012: waveform_sig_rx =244;
31013: waveform_sig_rx =461;
31014: waveform_sig_rx =336;
31015: waveform_sig_rx =260;
31016: waveform_sig_rx =278;
31017: waveform_sig_rx =502;
31018: waveform_sig_rx =160;
31019: waveform_sig_rx =233;
31020: waveform_sig_rx =511;
31021: waveform_sig_rx =147;
31022: waveform_sig_rx =185;
31023: waveform_sig_rx =451;
31024: waveform_sig_rx =232;
31025: waveform_sig_rx =104;
31026: waveform_sig_rx =378;
31027: waveform_sig_rx =278;
31028: waveform_sig_rx =100;
31029: waveform_sig_rx =241;
31030: waveform_sig_rx =346;
31031: waveform_sig_rx =95;
31032: waveform_sig_rx =217;
31033: waveform_sig_rx =163;
31034: waveform_sig_rx =241;
31035: waveform_sig_rx =146;
31036: waveform_sig_rx =217;
31037: waveform_sig_rx =165;
31038: waveform_sig_rx =1;
31039: waveform_sig_rx =421;
31040: waveform_sig_rx =-119;
31041: waveform_sig_rx =162;
31042: waveform_sig_rx =331;
31043: waveform_sig_rx =-183;
31044: waveform_sig_rx =226;
31045: waveform_sig_rx =274;
31046: waveform_sig_rx =-149;
31047: waveform_sig_rx =166;
31048: waveform_sig_rx =236;
31049: waveform_sig_rx =-100;
31050: waveform_sig_rx =110;
31051: waveform_sig_rx =147;
31052: waveform_sig_rx =25;
31053: waveform_sig_rx =-97;
31054: waveform_sig_rx =167;
31055: waveform_sig_rx =53;
31056: waveform_sig_rx =-122;
31057: waveform_sig_rx =25;
31058: waveform_sig_rx =185;
31059: waveform_sig_rx =-190;
31060: waveform_sig_rx =-2;
31061: waveform_sig_rx =166;
31062: waveform_sig_rx =-175;
31063: waveform_sig_rx =-80;
31064: waveform_sig_rx =133;
31065: waveform_sig_rx =-73;
31066: waveform_sig_rx =-160;
31067: waveform_sig_rx =53;
31068: waveform_sig_rx =-17;
31069: waveform_sig_rx =-191;
31070: waveform_sig_rx =-91;
31071: waveform_sig_rx =83;
31072: waveform_sig_rx =-241;
31073: waveform_sig_rx =-92;
31074: waveform_sig_rx =-102;
31075: waveform_sig_rx =-153;
31076: waveform_sig_rx =-140;
31077: waveform_sig_rx =-85;
31078: waveform_sig_rx =-225;
31079: waveform_sig_rx =-216;
31080: waveform_sig_rx =63;
31081: waveform_sig_rx =-445;
31082: waveform_sig_rx =-46;
31083: waveform_sig_rx =-78;
31084: waveform_sig_rx =-415;
31085: waveform_sig_rx =-48;
31086: waveform_sig_rx =-102;
31087: waveform_sig_rx =-388;
31088: waveform_sig_rx =-160;
31089: waveform_sig_rx =-81;
31090: waveform_sig_rx =-374;
31091: waveform_sig_rx =-238;
31092: waveform_sig_rx =-126;
31093: waveform_sig_rx =-280;
31094: waveform_sig_rx =-435;
31095: waveform_sig_rx =-91;
31096: waveform_sig_rx =-264;
31097: waveform_sig_rx =-450;
31098: waveform_sig_rx =-218;
31099: waveform_sig_rx =-159;
31100: waveform_sig_rx =-478;
31101: waveform_sig_rx =-249;
31102: waveform_sig_rx =-200;
31103: waveform_sig_rx =-428;
31104: waveform_sig_rx =-371;
31105: waveform_sig_rx =-220;
31106: waveform_sig_rx =-317;
31107: waveform_sig_rx =-493;
31108: waveform_sig_rx =-256;
31109: waveform_sig_rx =-272;
31110: waveform_sig_rx =-572;
31111: waveform_sig_rx =-351;
31112: waveform_sig_rx =-227;
31113: waveform_sig_rx =-609;
31114: waveform_sig_rx =-311;
31115: waveform_sig_rx =-448;
31116: waveform_sig_rx =-454;
31117: waveform_sig_rx =-373;
31118: waveform_sig_rx =-396;
31119: waveform_sig_rx =-495;
31120: waveform_sig_rx =-464;
31121: waveform_sig_rx =-303;
31122: waveform_sig_rx =-681;
31123: waveform_sig_rx =-348;
31124: waveform_sig_rx =-435;
31125: waveform_sig_rx =-648;
31126: waveform_sig_rx =-408;
31127: waveform_sig_rx =-372;
31128: waveform_sig_rx =-662;
31129: waveform_sig_rx =-505;
31130: waveform_sig_rx =-325;
31131: waveform_sig_rx =-696;
31132: waveform_sig_rx =-534;
31133: waveform_sig_rx =-381;
31134: waveform_sig_rx =-650;
31135: waveform_sig_rx =-709;
31136: waveform_sig_rx =-356;
31137: waveform_sig_rx =-629;
31138: waveform_sig_rx =-674;
31139: waveform_sig_rx =-515;
31140: waveform_sig_rx =-484;
31141: waveform_sig_rx =-738;
31142: waveform_sig_rx =-562;
31143: waveform_sig_rx =-469;
31144: waveform_sig_rx =-683;
31145: waveform_sig_rx =-695;
31146: waveform_sig_rx =-496;
31147: waveform_sig_rx =-600;
31148: waveform_sig_rx =-842;
31149: waveform_sig_rx =-482;
31150: waveform_sig_rx =-568;
31151: waveform_sig_rx =-863;
31152: waveform_sig_rx =-531;
31153: waveform_sig_rx =-532;
31154: waveform_sig_rx =-842;
31155: waveform_sig_rx =-545;
31156: waveform_sig_rx =-766;
31157: waveform_sig_rx =-649;
31158: waveform_sig_rx =-666;
31159: waveform_sig_rx =-716;
31160: waveform_sig_rx =-709;
31161: waveform_sig_rx =-758;
31162: waveform_sig_rx =-576;
31163: waveform_sig_rx =-886;
31164: waveform_sig_rx =-663;
31165: waveform_sig_rx =-608;
31166: waveform_sig_rx =-928;
31167: waveform_sig_rx =-705;
31168: waveform_sig_rx =-569;
31169: waveform_sig_rx =-1014;
31170: waveform_sig_rx =-720;
31171: waveform_sig_rx =-580;
31172: waveform_sig_rx =-1048;
31173: waveform_sig_rx =-736;
31174: waveform_sig_rx =-655;
31175: waveform_sig_rx =-913;
31176: waveform_sig_rx =-907;
31177: waveform_sig_rx =-644;
31178: waveform_sig_rx =-858;
31179: waveform_sig_rx =-918;
31180: waveform_sig_rx =-772;
31181: waveform_sig_rx =-738;
31182: waveform_sig_rx =-980;
31183: waveform_sig_rx =-839;
31184: waveform_sig_rx =-713;
31185: waveform_sig_rx =-927;
31186: waveform_sig_rx =-980;
31187: waveform_sig_rx =-648;
31188: waveform_sig_rx =-904;
31189: waveform_sig_rx =-1060;
31190: waveform_sig_rx =-635;
31191: waveform_sig_rx =-928;
31192: waveform_sig_rx =-1004;
31193: waveform_sig_rx =-780;
31194: waveform_sig_rx =-833;
31195: waveform_sig_rx =-992;
31196: waveform_sig_rx =-839;
31197: waveform_sig_rx =-965;
31198: waveform_sig_rx =-823;
31199: waveform_sig_rx =-965;
31200: waveform_sig_rx =-868;
31201: waveform_sig_rx =-963;
31202: waveform_sig_rx =-1006;
31203: waveform_sig_rx =-736;
31204: waveform_sig_rx =-1168;
31205: waveform_sig_rx =-887;
31206: waveform_sig_rx =-832;
31207: waveform_sig_rx =-1198;
31208: waveform_sig_rx =-877;
31209: waveform_sig_rx =-829;
31210: waveform_sig_rx =-1247;
31211: waveform_sig_rx =-891;
31212: waveform_sig_rx =-813;
31213: waveform_sig_rx =-1240;
31214: waveform_sig_rx =-906;
31215: waveform_sig_rx =-897;
31216: waveform_sig_rx =-1114;
31217: waveform_sig_rx =-1063;
31218: waveform_sig_rx =-854;
31219: waveform_sig_rx =-1052;
31220: waveform_sig_rx =-1078;
31221: waveform_sig_rx =-999;
31222: waveform_sig_rx =-888;
31223: waveform_sig_rx =-1176;
31224: waveform_sig_rx =-1017;
31225: waveform_sig_rx =-845;
31226: waveform_sig_rx =-1189;
31227: waveform_sig_rx =-1101;
31228: waveform_sig_rx =-825;
31229: waveform_sig_rx =-1160;
31230: waveform_sig_rx =-1141;
31231: waveform_sig_rx =-868;
31232: waveform_sig_rx =-1095;
31233: waveform_sig_rx =-1134;
31234: waveform_sig_rx =-1030;
31235: waveform_sig_rx =-940;
31236: waveform_sig_rx =-1171;
31237: waveform_sig_rx =-1050;
31238: waveform_sig_rx =-1085;
31239: waveform_sig_rx =-1051;
31240: waveform_sig_rx =-1116;
31241: waveform_sig_rx =-965;
31242: waveform_sig_rx =-1178;
31243: waveform_sig_rx =-1093;
31244: waveform_sig_rx =-920;
31245: waveform_sig_rx =-1343;
31246: waveform_sig_rx =-953;
31247: waveform_sig_rx =-1018;
31248: waveform_sig_rx =-1341;
31249: waveform_sig_rx =-965;
31250: waveform_sig_rx =-996;
31251: waveform_sig_rx =-1378;
31252: waveform_sig_rx =-955;
31253: waveform_sig_rx =-1007;
31254: waveform_sig_rx =-1348;
31255: waveform_sig_rx =-981;
31256: waveform_sig_rx =-1076;
31257: waveform_sig_rx =-1181;
31258: waveform_sig_rx =-1188;
31259: waveform_sig_rx =-997;
31260: waveform_sig_rx =-1113;
31261: waveform_sig_rx =-1264;
31262: waveform_sig_rx =-1051;
31263: waveform_sig_rx =-968;
31264: waveform_sig_rx =-1379;
31265: waveform_sig_rx =-1021;
31266: waveform_sig_rx =-1031;
31267: waveform_sig_rx =-1296;
31268: waveform_sig_rx =-1107;
31269: waveform_sig_rx =-1005;
31270: waveform_sig_rx =-1201;
31271: waveform_sig_rx =-1250;
31272: waveform_sig_rx =-1013;
31273: waveform_sig_rx =-1130;
31274: waveform_sig_rx =-1284;
31275: waveform_sig_rx =-1092;
31276: waveform_sig_rx =-1018;
31277: waveform_sig_rx =-1309;
31278: waveform_sig_rx =-1086;
31279: waveform_sig_rx =-1190;
31280: waveform_sig_rx =-1136;
31281: waveform_sig_rx =-1170;
31282: waveform_sig_rx =-1047;
31283: waveform_sig_rx =-1282;
31284: waveform_sig_rx =-1111;
31285: waveform_sig_rx =-1015;
31286: waveform_sig_rx =-1426;
31287: waveform_sig_rx =-959;
31288: waveform_sig_rx =-1125;
31289: waveform_sig_rx =-1380;
31290: waveform_sig_rx =-943;
31291: waveform_sig_rx =-1132;
31292: waveform_sig_rx =-1362;
31293: waveform_sig_rx =-1008;
31294: waveform_sig_rx =-1111;
31295: waveform_sig_rx =-1305;
31296: waveform_sig_rx =-1113;
31297: waveform_sig_rx =-1077;
31298: waveform_sig_rx =-1230;
31299: waveform_sig_rx =-1283;
31300: waveform_sig_rx =-961;
31301: waveform_sig_rx =-1217;
31302: waveform_sig_rx =-1291;
31303: waveform_sig_rx =-1037;
31304: waveform_sig_rx =-1085;
31305: waveform_sig_rx =-1364;
31306: waveform_sig_rx =-1045;
31307: waveform_sig_rx =-1090;
31308: waveform_sig_rx =-1283;
31309: waveform_sig_rx =-1164;
31310: waveform_sig_rx =-1046;
31311: waveform_sig_rx =-1212;
31312: waveform_sig_rx =-1256;
31313: waveform_sig_rx =-1008;
31314: waveform_sig_rx =-1117;
31315: waveform_sig_rx =-1314;
31316: waveform_sig_rx =-1059;
31317: waveform_sig_rx =-1024;
31318: waveform_sig_rx =-1354;
31319: waveform_sig_rx =-1018;
31320: waveform_sig_rx =-1209;
31321: waveform_sig_rx =-1128;
31322: waveform_sig_rx =-1145;
31323: waveform_sig_rx =-1101;
31324: waveform_sig_rx =-1273;
31325: waveform_sig_rx =-1063;
31326: waveform_sig_rx =-1064;
31327: waveform_sig_rx =-1372;
31328: waveform_sig_rx =-951;
31329: waveform_sig_rx =-1166;
31330: waveform_sig_rx =-1289;
31331: waveform_sig_rx =-989;
31332: waveform_sig_rx =-1101;
31333: waveform_sig_rx =-1303;
31334: waveform_sig_rx =-1038;
31335: waveform_sig_rx =-1019;
31336: waveform_sig_rx =-1300;
31337: waveform_sig_rx =-1081;
31338: waveform_sig_rx =-949;
31339: waveform_sig_rx =-1243;
31340: waveform_sig_rx =-1182;
31341: waveform_sig_rx =-905;
31342: waveform_sig_rx =-1234;
31343: waveform_sig_rx =-1181;
31344: waveform_sig_rx =-995;
31345: waveform_sig_rx =-1066;
31346: waveform_sig_rx =-1268;
31347: waveform_sig_rx =-1010;
31348: waveform_sig_rx =-1019;
31349: waveform_sig_rx =-1207;
31350: waveform_sig_rx =-1110;
31351: waveform_sig_rx =-945;
31352: waveform_sig_rx =-1123;
31353: waveform_sig_rx =-1223;
31354: waveform_sig_rx =-905;
31355: waveform_sig_rx =-1062;
31356: waveform_sig_rx =-1284;
31357: waveform_sig_rx =-903;
31358: waveform_sig_rx =-1015;
31359: waveform_sig_rx =-1250;
31360: waveform_sig_rx =-883;
31361: waveform_sig_rx =-1227;
31362: waveform_sig_rx =-949;
31363: waveform_sig_rx =-1097;
31364: waveform_sig_rx =-1012;
31365: waveform_sig_rx =-1112;
31366: waveform_sig_rx =-1008;
31367: waveform_sig_rx =-942;
31368: waveform_sig_rx =-1228;
31369: waveform_sig_rx =-905;
31370: waveform_sig_rx =-997;
31371: waveform_sig_rx =-1217;
31372: waveform_sig_rx =-865;
31373: waveform_sig_rx =-962;
31374: waveform_sig_rx =-1227;
31375: waveform_sig_rx =-880;
31376: waveform_sig_rx =-920;
31377: waveform_sig_rx =-1197;
31378: waveform_sig_rx =-944;
31379: waveform_sig_rx =-863;
31380: waveform_sig_rx =-1169;
31381: waveform_sig_rx =-1033;
31382: waveform_sig_rx =-789;
31383: waveform_sig_rx =-1141;
31384: waveform_sig_rx =-994;
31385: waveform_sig_rx =-912;
31386: waveform_sig_rx =-922;
31387: waveform_sig_rx =-1069;
31388: waveform_sig_rx =-926;
31389: waveform_sig_rx =-817;
31390: waveform_sig_rx =-1082;
31391: waveform_sig_rx =-975;
31392: waveform_sig_rx =-734;
31393: waveform_sig_rx =-1061;
31394: waveform_sig_rx =-1033;
31395: waveform_sig_rx =-710;
31396: waveform_sig_rx =-986;
31397: waveform_sig_rx =-1043;
31398: waveform_sig_rx =-765;
31399: waveform_sig_rx =-892;
31400: waveform_sig_rx =-1020;
31401: waveform_sig_rx =-790;
31402: waveform_sig_rx =-1026;
31403: waveform_sig_rx =-772;
31404: waveform_sig_rx =-984;
31405: waveform_sig_rx =-808;
31406: waveform_sig_rx =-993;
31407: waveform_sig_rx =-854;
31408: waveform_sig_rx =-767;
31409: waveform_sig_rx =-1081;
31410: waveform_sig_rx =-711;
31411: waveform_sig_rx =-839;
31412: waveform_sig_rx =-1068;
31413: waveform_sig_rx =-687;
31414: waveform_sig_rx =-785;
31415: waveform_sig_rx =-1091;
31416: waveform_sig_rx =-672;
31417: waveform_sig_rx =-745;
31418: waveform_sig_rx =-1060;
31419: waveform_sig_rx =-689;
31420: waveform_sig_rx =-700;
31421: waveform_sig_rx =-996;
31422: waveform_sig_rx =-767;
31423: waveform_sig_rx =-660;
31424: waveform_sig_rx =-883;
31425: waveform_sig_rx =-790;
31426: waveform_sig_rx =-754;
31427: waveform_sig_rx =-641;
31428: waveform_sig_rx =-953;
31429: waveform_sig_rx =-688;
31430: waveform_sig_rx =-600;
31431: waveform_sig_rx =-964;
31432: waveform_sig_rx =-704;
31433: waveform_sig_rx =-569;
31434: waveform_sig_rx =-877;
31435: waveform_sig_rx =-762;
31436: waveform_sig_rx =-598;
31437: waveform_sig_rx =-771;
31438: waveform_sig_rx =-829;
31439: waveform_sig_rx =-582;
31440: waveform_sig_rx =-673;
31441: waveform_sig_rx =-815;
31442: waveform_sig_rx =-574;
31443: waveform_sig_rx =-801;
31444: waveform_sig_rx =-538;
31445: waveform_sig_rx =-758;
31446: waveform_sig_rx =-541;
31447: waveform_sig_rx =-782;
31448: waveform_sig_rx =-600;
31449: waveform_sig_rx =-510;
31450: waveform_sig_rx =-888;
31451: waveform_sig_rx =-445;
31452: waveform_sig_rx =-610;
31453: waveform_sig_rx =-865;
31454: waveform_sig_rx =-360;
31455: waveform_sig_rx =-619;
31456: waveform_sig_rx =-831;
31457: waveform_sig_rx =-370;
31458: waveform_sig_rx =-615;
31459: waveform_sig_rx =-728;
31460: waveform_sig_rx =-444;
31461: waveform_sig_rx =-520;
31462: waveform_sig_rx =-687;
31463: waveform_sig_rx =-572;
31464: waveform_sig_rx =-438;
31465: waveform_sig_rx =-590;
31466: waveform_sig_rx =-619;
31467: waveform_sig_rx =-451;
31468: waveform_sig_rx =-425;
31469: waveform_sig_rx =-749;
31470: waveform_sig_rx =-353;
31471: waveform_sig_rx =-427;
31472: waveform_sig_rx =-677;
31473: waveform_sig_rx =-412;
31474: waveform_sig_rx =-366;
31475: waveform_sig_rx =-592;
31476: waveform_sig_rx =-511;
31477: waveform_sig_rx =-333;
31478: waveform_sig_rx =-494;
31479: waveform_sig_rx =-581;
31480: waveform_sig_rx =-327;
31481: waveform_sig_rx =-403;
31482: waveform_sig_rx =-550;
31483: waveform_sig_rx =-354;
31484: waveform_sig_rx =-507;
31485: waveform_sig_rx =-335;
31486: waveform_sig_rx =-500;
31487: waveform_sig_rx =-266;
31488: waveform_sig_rx =-589;
31489: waveform_sig_rx =-284;
31490: waveform_sig_rx =-307;
31491: waveform_sig_rx =-629;
31492: waveform_sig_rx =-91;
31493: waveform_sig_rx =-433;
31494: waveform_sig_rx =-548;
31495: waveform_sig_rx =-84;
31496: waveform_sig_rx =-425;
31497: waveform_sig_rx =-470;
31498: waveform_sig_rx =-139;
31499: waveform_sig_rx =-331;
31500: waveform_sig_rx =-415;
31501: waveform_sig_rx =-233;
31502: waveform_sig_rx =-211;
31503: waveform_sig_rx =-435;
31504: waveform_sig_rx =-301;
31505: waveform_sig_rx =-107;
31506: waveform_sig_rx =-365;
31507: waveform_sig_rx =-340;
31508: waveform_sig_rx =-143;
31509: waveform_sig_rx =-182;
31510: waveform_sig_rx =-458;
31511: waveform_sig_rx =-54;
31512: waveform_sig_rx =-163;
31513: waveform_sig_rx =-401;
31514: waveform_sig_rx =-118;
31515: waveform_sig_rx =-116;
31516: waveform_sig_rx =-291;
31517: waveform_sig_rx =-247;
31518: waveform_sig_rx =-70;
31519: waveform_sig_rx =-207;
31520: waveform_sig_rx =-347;
31521: waveform_sig_rx =-22;
31522: waveform_sig_rx =-120;
31523: waveform_sig_rx =-322;
31524: waveform_sig_rx =-24;
31525: waveform_sig_rx =-242;
31526: waveform_sig_rx =-55;
31527: waveform_sig_rx =-159;
31528: waveform_sig_rx =-34;
31529: waveform_sig_rx =-302;
31530: waveform_sig_rx =55;
31531: waveform_sig_rx =-91;
31532: waveform_sig_rx =-282;
31533: waveform_sig_rx =163;
31534: waveform_sig_rx =-171;
31535: waveform_sig_rx =-167;
31536: waveform_sig_rx =142;
31537: waveform_sig_rx =-92;
31538: waveform_sig_rx =-173;
31539: waveform_sig_rx =126;
31540: waveform_sig_rx =-12;
31541: waveform_sig_rx =-154;
31542: waveform_sig_rx =73;
31543: waveform_sig_rx =104;
31544: waveform_sig_rx =-164;
31545: waveform_sig_rx =5;
31546: waveform_sig_rx =195;
31547: waveform_sig_rx =-95;
31548: waveform_sig_rx =-49;
31549: waveform_sig_rx =178;
31550: waveform_sig_rx =45;
31551: waveform_sig_rx =-129;
31552: waveform_sig_rx =201;
31553: waveform_sig_rx =80;
31554: waveform_sig_rx =-68;
31555: waveform_sig_rx =109;
31556: waveform_sig_rx =197;
31557: waveform_sig_rx =5;
31558: waveform_sig_rx =9;
31559: waveform_sig_rx =276;
31560: waveform_sig_rx =55;
31561: waveform_sig_rx =-41;
31562: waveform_sig_rx =334;
31563: waveform_sig_rx =136;
31564: waveform_sig_rx =6;
31565: waveform_sig_rx =287;
31566: waveform_sig_rx =22;
31567: waveform_sig_rx =282;
31568: waveform_sig_rx =124;
31569: waveform_sig_rx =241;
31570: waveform_sig_rx =57;
31571: waveform_sig_rx =338;
31572: waveform_sig_rx =178;
31573: waveform_sig_rx =71;
31574: waveform_sig_rx =405;
31575: waveform_sig_rx =141;
31576: waveform_sig_rx =107;
31577: waveform_sig_rx =387;
31578: waveform_sig_rx =233;
31579: waveform_sig_rx =59;
31580: waveform_sig_rx =425;
31581: waveform_sig_rx =299;
31582: waveform_sig_rx =86;
31583: waveform_sig_rx =392;
31584: waveform_sig_rx =391;
31585: waveform_sig_rx =75;
31586: waveform_sig_rx =339;
31587: waveform_sig_rx =438;
31588: waveform_sig_rx =178;
31589: waveform_sig_rx =287;
31590: waveform_sig_rx =433;
31591: waveform_sig_rx =321;
31592: waveform_sig_rx =206;
31593: waveform_sig_rx =482;
31594: waveform_sig_rx =378;
31595: waveform_sig_rx =242;
31596: waveform_sig_rx =381;
31597: waveform_sig_rx =525;
31598: waveform_sig_rx =239;
31599: waveform_sig_rx =309;
31600: waveform_sig_rx =606;
31601: waveform_sig_rx =282;
31602: waveform_sig_rx =296;
31603: waveform_sig_rx =606;
31604: waveform_sig_rx =372;
31605: waveform_sig_rx =342;
31606: waveform_sig_rx =539;
31607: waveform_sig_rx =318;
31608: waveform_sig_rx =570;
31609: waveform_sig_rx =363;
31610: waveform_sig_rx =542;
31611: waveform_sig_rx =337;
31612: waveform_sig_rx =574;
31613: waveform_sig_rx =477;
31614: waveform_sig_rx =350;
31615: waveform_sig_rx =661;
31616: waveform_sig_rx =469;
31617: waveform_sig_rx =356;
31618: waveform_sig_rx =721;
31619: waveform_sig_rx =513;
31620: waveform_sig_rx =306;
31621: waveform_sig_rx =785;
31622: waveform_sig_rx =516;
31623: waveform_sig_rx =379;
31624: waveform_sig_rx =704;
31625: waveform_sig_rx =613;
31626: waveform_sig_rx =391;
31627: waveform_sig_rx =625;
31628: waveform_sig_rx =689;
31629: waveform_sig_rx =466;
31630: waveform_sig_rx =545;
31631: waveform_sig_rx =715;
31632: waveform_sig_rx =593;
31633: waveform_sig_rx =479;
31634: waveform_sig_rx =733;
31635: waveform_sig_rx =668;
31636: waveform_sig_rx =475;
31637: waveform_sig_rx =655;
31638: waveform_sig_rx =818;
31639: waveform_sig_rx =447;
31640: waveform_sig_rx =639;
31641: waveform_sig_rx =862;
31642: waveform_sig_rx =497;
31643: waveform_sig_rx =648;
31644: waveform_sig_rx =806;
31645: waveform_sig_rx =629;
31646: waveform_sig_rx =661;
31647: waveform_sig_rx =710;
31648: waveform_sig_rx =650;
31649: waveform_sig_rx =791;
31650: waveform_sig_rx =614;
31651: waveform_sig_rx =840;
31652: waveform_sig_rx =540;
31653: waveform_sig_rx =882;
31654: waveform_sig_rx =732;
31655: waveform_sig_rx =552;
31656: waveform_sig_rx =951;
31657: waveform_sig_rx =673;
31658: waveform_sig_rx =606;
31659: waveform_sig_rx =992;
31660: waveform_sig_rx =711;
31661: waveform_sig_rx =569;
31662: waveform_sig_rx =1014;
31663: waveform_sig_rx =717;
31664: waveform_sig_rx =622;
31665: waveform_sig_rx =967;
31666: waveform_sig_rx =807;
31667: waveform_sig_rx =635;
31668: waveform_sig_rx =884;
31669: waveform_sig_rx =884;
31670: waveform_sig_rx =744;
31671: waveform_sig_rx =772;
31672: waveform_sig_rx =953;
31673: waveform_sig_rx =862;
31674: waveform_sig_rx =649;
31675: waveform_sig_rx =1019;
31676: waveform_sig_rx =871;
31677: waveform_sig_rx =673;
31678: waveform_sig_rx =957;
31679: waveform_sig_rx =969;
31680: waveform_sig_rx =675;
31681: waveform_sig_rx =902;
31682: waveform_sig_rx =995;
31683: waveform_sig_rx =775;
31684: waveform_sig_rx =844;
31685: waveform_sig_rx =1005;
31686: waveform_sig_rx =901;
31687: waveform_sig_rx =820;
31688: waveform_sig_rx =954;
31689: waveform_sig_rx =883;
31690: waveform_sig_rx =966;
31691: waveform_sig_rx =865;
31692: waveform_sig_rx =1019;
31693: waveform_sig_rx =725;
31694: waveform_sig_rx =1134;
31695: waveform_sig_rx =877;
31696: waveform_sig_rx =796;
31697: waveform_sig_rx =1171;
31698: waveform_sig_rx =833;
31699: waveform_sig_rx =828;
31700: waveform_sig_rx =1178;
31701: waveform_sig_rx =862;
31702: waveform_sig_rx =774;
31703: waveform_sig_rx =1232;
31704: waveform_sig_rx =847;
31705: waveform_sig_rx =857;
31706: waveform_sig_rx =1143;
31707: waveform_sig_rx =946;
31708: waveform_sig_rx =870;
31709: waveform_sig_rx =1009;
31710: waveform_sig_rx =1093;
31711: waveform_sig_rx =932;
31712: waveform_sig_rx =875;
31713: waveform_sig_rx =1211;
31714: waveform_sig_rx =959;
31715: waveform_sig_rx =849;
31716: waveform_sig_rx =1238;
31717: waveform_sig_rx =945;
31718: waveform_sig_rx =904;
31719: waveform_sig_rx =1105;
31720: waveform_sig_rx =1087;
31721: waveform_sig_rx =907;
31722: waveform_sig_rx =1008;
31723: waveform_sig_rx =1202;
31724: waveform_sig_rx =926;
31725: waveform_sig_rx =963;
31726: waveform_sig_rx =1230;
31727: waveform_sig_rx =996;
31728: waveform_sig_rx =965;
31729: waveform_sig_rx =1108;
31730: waveform_sig_rx =1002;
31731: waveform_sig_rx =1114;
31732: waveform_sig_rx =1008;
31733: waveform_sig_rx =1165;
31734: waveform_sig_rx =861;
31735: waveform_sig_rx =1297;
31736: waveform_sig_rx =990;
31737: waveform_sig_rx =956;
31738: waveform_sig_rx =1311;
31739: waveform_sig_rx =906;
31740: waveform_sig_rx =1012;
31741: waveform_sig_rx =1327;
31742: waveform_sig_rx =937;
31743: waveform_sig_rx =999;
31744: waveform_sig_rx =1302;
31745: waveform_sig_rx =977;
31746: waveform_sig_rx =1036;
31747: waveform_sig_rx =1167;
31748: waveform_sig_rx =1156;
31749: waveform_sig_rx =934;
31750: waveform_sig_rx =1137;
31751: waveform_sig_rx =1257;
31752: waveform_sig_rx =943;
31753: waveform_sig_rx =1085;
31754: waveform_sig_rx =1297;
31755: waveform_sig_rx =1001;
31756: waveform_sig_rx =1047;
31757: waveform_sig_rx =1268;
31758: waveform_sig_rx =1088;
31759: waveform_sig_rx =1022;
31760: waveform_sig_rx =1173;
31761: waveform_sig_rx =1240;
31762: waveform_sig_rx =954;
31763: waveform_sig_rx =1135;
31764: waveform_sig_rx =1280;
31765: waveform_sig_rx =1013;
31766: waveform_sig_rx =1067;
31767: waveform_sig_rx =1315;
31768: waveform_sig_rx =1078;
31769: waveform_sig_rx =1074;
31770: waveform_sig_rx =1220;
31771: waveform_sig_rx =1062;
31772: waveform_sig_rx =1203;
31773: waveform_sig_rx =1129;
31774: waveform_sig_rx =1180;
31775: waveform_sig_rx =977;
31776: waveform_sig_rx =1363;
31777: waveform_sig_rx =998;
31778: waveform_sig_rx =1097;
31779: waveform_sig_rx =1324;
31780: waveform_sig_rx =984;
31781: waveform_sig_rx =1117;
31782: waveform_sig_rx =1310;
31783: waveform_sig_rx =1067;
31784: waveform_sig_rx =1019;
31785: waveform_sig_rx =1385;
31786: waveform_sig_rx =1070;
31787: waveform_sig_rx =1036;
31788: waveform_sig_rx =1295;
31789: waveform_sig_rx =1201;
31790: waveform_sig_rx =956;
31791: waveform_sig_rx =1267;
31792: waveform_sig_rx =1222;
31793: waveform_sig_rx =1014;
31794: waveform_sig_rx =1161;
31795: waveform_sig_rx =1291;
31796: waveform_sig_rx =1072;
31797: waveform_sig_rx =1081;
31798: waveform_sig_rx =1309;
31799: waveform_sig_rx =1131;
31800: waveform_sig_rx =1052;
31801: waveform_sig_rx =1244;
31802: waveform_sig_rx =1273;
31803: waveform_sig_rx =986;
31804: waveform_sig_rx =1167;
31805: waveform_sig_rx =1335;
31806: waveform_sig_rx =1011;
31807: waveform_sig_rx =1092;
31808: waveform_sig_rx =1360;
31809: waveform_sig_rx =1014;
31810: waveform_sig_rx =1137;
31811: waveform_sig_rx =1230;
31812: waveform_sig_rx =1030;
31813: waveform_sig_rx =1273;
31814: waveform_sig_rx =1086;
31815: waveform_sig_rx =1203;
31816: waveform_sig_rx =1036;
31817: waveform_sig_rx =1330;
31818: waveform_sig_rx =1046;
31819: waveform_sig_rx =1083;
31820: waveform_sig_rx =1318;
31821: waveform_sig_rx =1050;
31822: waveform_sig_rx =1061;
31823: waveform_sig_rx =1340;
31824: waveform_sig_rx =1052;
31825: waveform_sig_rx =994;
31826: waveform_sig_rx =1392;
31827: waveform_sig_rx =1011;
31828: waveform_sig_rx =1039;
31829: waveform_sig_rx =1294;
31830: waveform_sig_rx =1125;
31831: waveform_sig_rx =929;
31832: waveform_sig_rx =1254;
31833: waveform_sig_rx =1173;
31834: waveform_sig_rx =999;
31835: waveform_sig_rx =1131;
31836: waveform_sig_rx =1236;
31837: waveform_sig_rx =1059;
31838: waveform_sig_rx =1028;
31839: waveform_sig_rx =1266;
31840: waveform_sig_rx =1101;
31841: waveform_sig_rx =968;
31842: waveform_sig_rx =1201;
31843: waveform_sig_rx =1206;
31844: waveform_sig_rx =881;
31845: waveform_sig_rx =1159;
31846: waveform_sig_rx =1227;
31847: waveform_sig_rx =920;
31848: waveform_sig_rx =1093;
31849: waveform_sig_rx =1257;
31850: waveform_sig_rx =978;
31851: waveform_sig_rx =1131;
31852: waveform_sig_rx =1088;
31853: waveform_sig_rx =1051;
31854: waveform_sig_rx =1165;
31855: waveform_sig_rx =976;
31856: waveform_sig_rx =1166;
31857: waveform_sig_rx =890;
31858: waveform_sig_rx =1254;
31859: waveform_sig_rx =962;
31860: waveform_sig_rx =971;
31861: waveform_sig_rx =1259;
31862: waveform_sig_rx =905;
31863: waveform_sig_rx =973;
31864: waveform_sig_rx =1284;
31865: waveform_sig_rx =887;
31866: waveform_sig_rx =940;
31867: waveform_sig_rx =1295;
31868: waveform_sig_rx =877;
31869: waveform_sig_rx =962;
31870: waveform_sig_rx =1210;
31871: waveform_sig_rx =979;
31872: waveform_sig_rx =865;
31873: waveform_sig_rx =1180;
31874: waveform_sig_rx =1025;
31875: waveform_sig_rx =945;
31876: waveform_sig_rx =975;
31877: waveform_sig_rx =1144;
31878: waveform_sig_rx =963;
31879: waveform_sig_rx =861;
31880: waveform_sig_rx =1203;
31881: waveform_sig_rx =947;
31882: waveform_sig_rx =823;
31883: waveform_sig_rx =1155;
31884: waveform_sig_rx =1009;
31885: waveform_sig_rx =807;
31886: waveform_sig_rx =1083;
31887: waveform_sig_rx =1067;
31888: waveform_sig_rx =835;
31889: waveform_sig_rx =962;
31890: waveform_sig_rx =1130;
31891: waveform_sig_rx =846;
31892: waveform_sig_rx =967;
31893: waveform_sig_rx =947;
31894: waveform_sig_rx =939;
31895: waveform_sig_rx =996;
31896: waveform_sig_rx =880;
31897: waveform_sig_rx =1025;
31898: waveform_sig_rx =724;
31899: waveform_sig_rx =1139;
31900: waveform_sig_rx =797;
31901: waveform_sig_rx =810;
31902: waveform_sig_rx =1146;
31903: waveform_sig_rx =676;
31904: waveform_sig_rx =853;
31905: waveform_sig_rx =1149;
31906: waveform_sig_rx =654;
31907: waveform_sig_rx =861;
31908: waveform_sig_rx =1080;
31909: waveform_sig_rx =705;
31910: waveform_sig_rx =873;
31911: waveform_sig_rx =962;
31912: waveform_sig_rx =844;
31913: waveform_sig_rx =705;
31914: waveform_sig_rx =952;
31915: waveform_sig_rx =876;
31916: waveform_sig_rx =730;
31917: waveform_sig_rx =791;
31918: waveform_sig_rx =997;
31919: waveform_sig_rx =718;
31920: waveform_sig_rx =698;
31921: waveform_sig_rx =1033;
31922: waveform_sig_rx =717;
31923: waveform_sig_rx =678;
31924: waveform_sig_rx =955;
31925: waveform_sig_rx =794;
31926: waveform_sig_rx =658;
31927: waveform_sig_rx =840;
31928: waveform_sig_rx =843;
31929: waveform_sig_rx =661;
31930: waveform_sig_rx =715;
31931: waveform_sig_rx =932;
31932: waveform_sig_rx =647;
31933: waveform_sig_rx =735;
31934: waveform_sig_rx =758;
31935: waveform_sig_rx =692;
31936: waveform_sig_rx =754;
31937: waveform_sig_rx =708;
31938: waveform_sig_rx =757;
31939: waveform_sig_rx =533;
31940: waveform_sig_rx =966;
31941: waveform_sig_rx =488;
31942: waveform_sig_rx =659;
31943: waveform_sig_rx =926;
31944: waveform_sig_rx =416;
31945: waveform_sig_rx =735;
31946: waveform_sig_rx =860;
31947: waveform_sig_rx =425;
31948: waveform_sig_rx =683;
31949: waveform_sig_rx =800;
31950: waveform_sig_rx =511;
31951: waveform_sig_rx =609;
31952: waveform_sig_rx =712;
31953: waveform_sig_rx =648;
31954: waveform_sig_rx =424;
31955: waveform_sig_rx =748;
31956: waveform_sig_rx =650;
31957: waveform_sig_rx =497;
31958: waveform_sig_rx =590;
31959: waveform_sig_rx =747;
31960: waveform_sig_rx =466;
31961: waveform_sig_rx =515;
31962: waveform_sig_rx =788;
31963: waveform_sig_rx =453;
31964: waveform_sig_rx =468;
31965: waveform_sig_rx =704;
31966: waveform_sig_rx =531;
31967: waveform_sig_rx =460;
31968: waveform_sig_rx =574;
31969: waveform_sig_rx =627;
31970: waveform_sig_rx =409;
31971: waveform_sig_rx =442;
31972: waveform_sig_rx =733;
31973: waveform_sig_rx =321;
31974: waveform_sig_rx =502;
31975: waveform_sig_rx =531;
31976: waveform_sig_rx =390;
31977: waveform_sig_rx =543;
31978: waveform_sig_rx =455;
31979: waveform_sig_rx =465;
31980: waveform_sig_rx =351;
31981: waveform_sig_rx =671;
31982: waveform_sig_rx =235;
31983: waveform_sig_rx =469;
31984: waveform_sig_rx =595;
31985: waveform_sig_rx =196;
31986: waveform_sig_rx =471;
31987: waveform_sig_rx =571;
31988: waveform_sig_rx =210;
31989: waveform_sig_rx =407;
31990: waveform_sig_rx =542;
31991: waveform_sig_rx =249;
31992: waveform_sig_rx =350;
31993: waveform_sig_rx =472;
31994: waveform_sig_rx =391;
31995: waveform_sig_rx =133;
31996: waveform_sig_rx =510;
31997: waveform_sig_rx =367;
31998: waveform_sig_rx =170;
31999: waveform_sig_rx =363;
32000: waveform_sig_rx =438;
32001: waveform_sig_rx =169;
32002: waveform_sig_rx =284;
32003: waveform_sig_rx =428;
32004: waveform_sig_rx =191;
32005: waveform_sig_rx =209;
32006: waveform_sig_rx =386;
32007: waveform_sig_rx =300;
32008: waveform_sig_rx =84;
32009: waveform_sig_rx =293;
32010: waveform_sig_rx =364;
32011: waveform_sig_rx =40;
32012: waveform_sig_rx =220;
32013: waveform_sig_rx =411;
32014: waveform_sig_rx =5;
32015: waveform_sig_rx =291;
32016: waveform_sig_rx =175;
32017: waveform_sig_rx =133;
32018: waveform_sig_rx =249;
32019: waveform_sig_rx =130;
32020: waveform_sig_rx =177;
32021: waveform_sig_rx =66;
32022: waveform_sig_rx =344;
32023: waveform_sig_rx =-51;
32024: waveform_sig_rx =166;
32025: waveform_sig_rx =267;
32026: waveform_sig_rx =-69;
32027: waveform_sig_rx =153;
32028: waveform_sig_rx =250;
32029: waveform_sig_rx =-73;
32030: waveform_sig_rx =65;
32031: waveform_sig_rx =269;
32032: waveform_sig_rx =-76;
32033: waveform_sig_rx =-1;
32034: waveform_sig_rx =209;
32035: waveform_sig_rx =16;
32036: waveform_sig_rx =-153;
32037: waveform_sig_rx =240;
32038: waveform_sig_rx =5;
32039: waveform_sig_rx =-81;
32040: waveform_sig_rx =61;
32041: waveform_sig_rx =102;
32042: waveform_sig_rx =-101;
32043: waveform_sig_rx =-26;
32044: waveform_sig_rx =144;
32045: waveform_sig_rx =-84;
32046: waveform_sig_rx =-132;
32047: waveform_sig_rx =98;
32048: waveform_sig_rx =-16;
32049: waveform_sig_rx =-252;
32050: waveform_sig_rx =58;
32051: waveform_sig_rx =32;
32052: waveform_sig_rx =-288;
32053: waveform_sig_rx =-38;
32054: waveform_sig_rx =62;
32055: waveform_sig_rx =-292;
32056: waveform_sig_rx =-14;
32057: waveform_sig_rx =-173;
32058: waveform_sig_rx =-118;
32059: waveform_sig_rx =-80;
32060: waveform_sig_rx =-169;
32061: waveform_sig_rx =-102;
32062: waveform_sig_rx =-259;
32063: waveform_sig_rx =38;
32064: waveform_sig_rx =-311;
32065: waveform_sig_rx =-147;
32066: waveform_sig_rx =-25;
32067: waveform_sig_rx =-360;
32068: waveform_sig_rx =-174;
32069: waveform_sig_rx =0;
32070: waveform_sig_rx =-412;
32071: waveform_sig_rx =-225;
32072: waveform_sig_rx =9;
32073: waveform_sig_rx =-445;
32074: waveform_sig_rx =-235;
32075: waveform_sig_rx =-76;
32076: waveform_sig_rx =-345;
32077: waveform_sig_rx =-381;
32078: waveform_sig_rx =-110;
32079: waveform_sig_rx =-315;
32080: waveform_sig_rx =-360;
32081: waveform_sig_rx =-314;
32082: waveform_sig_rx =-163;
32083: waveform_sig_rx =-442;
32084: waveform_sig_rx =-359;
32085: waveform_sig_rx =-157;
32086: waveform_sig_rx =-417;
32087: waveform_sig_rx =-440;
32088: waveform_sig_rx =-183;
32089: waveform_sig_rx =-340;
32090: waveform_sig_rx =-542;
32091: waveform_sig_rx =-199;
32092: waveform_sig_rx =-312;
32093: waveform_sig_rx =-543;
32094: waveform_sig_rx =-293;
32095: waveform_sig_rx =-304;
32096: waveform_sig_rx =-522;
32097: waveform_sig_rx =-338;
32098: waveform_sig_rx =-508;
32099: waveform_sig_rx =-342;
32100: waveform_sig_rx =-456;
32101: waveform_sig_rx =-427;
32102: waveform_sig_rx =-419;
32103: waveform_sig_rx =-584;
32104: waveform_sig_rx =-227;
32105: waveform_sig_rx =-682;
32106: waveform_sig_rx =-463;
32107: waveform_sig_rx =-291;
32108: waveform_sig_rx =-718;
32109: waveform_sig_rx =-413;
32110: waveform_sig_rx =-320;
32111: waveform_sig_rx =-735;
32112: waveform_sig_rx =-473;
32113: waveform_sig_rx =-334;
32114: waveform_sig_rx =-730;
32115: waveform_sig_rx =-509;
32116: waveform_sig_rx =-393;
32117: waveform_sig_rx =-616;
32118: waveform_sig_rx =-655;
32119: waveform_sig_rx =-385;
32120: waveform_sig_rx =-592;
32121: waveform_sig_rx =-637;
32122: waveform_sig_rx =-592;
32123: waveform_sig_rx =-422;
32124: waveform_sig_rx =-736;
32125: waveform_sig_rx =-638;
32126: waveform_sig_rx =-401;
32127: waveform_sig_rx =-752;
32128: waveform_sig_rx =-689;
32129: waveform_sig_rx =-422;
32130: waveform_sig_rx =-684;
32131: waveform_sig_rx =-756;
32132: waveform_sig_rx =-495;
32133: waveform_sig_rx =-623;
32134: waveform_sig_rx =-755;
32135: waveform_sig_rx =-633;
32136: waveform_sig_rx =-510;
32137: waveform_sig_rx =-793;
32138: waveform_sig_rx =-646;
32139: waveform_sig_rx =-683;
32140: waveform_sig_rx =-657;
32141: waveform_sig_rx =-738;
32142: waveform_sig_rx =-646;
32143: waveform_sig_rx =-771;
32144: waveform_sig_rx =-788;
32145: waveform_sig_rx =-494;
32146: waveform_sig_rx =-973;
32147: waveform_sig_rx =-627;
32148: waveform_sig_rx =-592;
32149: waveform_sig_rx =-961;
32150: waveform_sig_rx =-651;
32151: waveform_sig_rx =-585;
32152: waveform_sig_rx =-1001;
32153: waveform_sig_rx =-690;
32154: waveform_sig_rx =-598;
32155: waveform_sig_rx =-1010;
32156: waveform_sig_rx =-707;
32157: waveform_sig_rx =-707;
32158: waveform_sig_rx =-852;
32159: waveform_sig_rx =-882;
32160: waveform_sig_rx =-706;
32161: waveform_sig_rx =-775;
32162: waveform_sig_rx =-959;
32163: waveform_sig_rx =-804;
32164: waveform_sig_rx =-628;
32165: waveform_sig_rx =-1072;
32166: waveform_sig_rx =-785;
32167: waveform_sig_rx =-685;
32168: waveform_sig_rx =-989;
32169: waveform_sig_rx =-849;
32170: waveform_sig_rx =-748;
32171: waveform_sig_rx =-856;
32172: waveform_sig_rx =-1000;
32173: waveform_sig_rx =-745;
32174: waveform_sig_rx =-796;
32175: waveform_sig_rx =-1051;
32176: waveform_sig_rx =-841;
32177: waveform_sig_rx =-731;
32178: waveform_sig_rx =-1056;
32179: waveform_sig_rx =-826;
32180: waveform_sig_rx =-920;
32181: waveform_sig_rx =-880;
32182: waveform_sig_rx =-917;
32183: waveform_sig_rx =-850;
32184: waveform_sig_rx =-1001;
32185: waveform_sig_rx =-970;
32186: waveform_sig_rx =-744;
32187: waveform_sig_rx =-1189;
32188: waveform_sig_rx =-822;
32189: waveform_sig_rx =-855;
32190: waveform_sig_rx =-1177;
32191: waveform_sig_rx =-823;
32192: waveform_sig_rx =-858;
32193: waveform_sig_rx =-1189;
32194: waveform_sig_rx =-889;
32195: waveform_sig_rx =-864;
32196: waveform_sig_rx =-1140;
32197: waveform_sig_rx =-951;
32198: waveform_sig_rx =-899;
32199: waveform_sig_rx =-999;
32200: waveform_sig_rx =-1170;
32201: waveform_sig_rx =-826;
32202: waveform_sig_rx =-997;
32203: waveform_sig_rx =-1201;
32204: waveform_sig_rx =-895;
32205: waveform_sig_rx =-926;
32206: waveform_sig_rx =-1222;
32207: waveform_sig_rx =-930;
32208: waveform_sig_rx =-964;
32209: waveform_sig_rx =-1113;
32210: waveform_sig_rx =-1096;
32211: waveform_sig_rx =-923;
32212: waveform_sig_rx =-1028;
32213: waveform_sig_rx =-1219;
32214: waveform_sig_rx =-873;
32215: waveform_sig_rx =-1015;
32216: waveform_sig_rx =-1226;
32217: waveform_sig_rx =-963;
32218: waveform_sig_rx =-932;
32219: waveform_sig_rx =-1206;
32220: waveform_sig_rx =-987;
32221: waveform_sig_rx =-1108;
32222: waveform_sig_rx =-1051;
32223: waveform_sig_rx =-1097;
32224: waveform_sig_rx =-1011;
32225: waveform_sig_rx =-1180;
32226: waveform_sig_rx =-1055;
32227: waveform_sig_rx =-946;
32228: waveform_sig_rx =-1327;
32229: waveform_sig_rx =-914;
32230: waveform_sig_rx =-1079;
32231: waveform_sig_rx =-1267;
32232: waveform_sig_rx =-1005;
32233: waveform_sig_rx =-1038;
32234: waveform_sig_rx =-1253;
32235: waveform_sig_rx =-1113;
32236: waveform_sig_rx =-918;
32237: waveform_sig_rx =-1296;
32238: waveform_sig_rx =-1103;
32239: waveform_sig_rx =-933;
32240: waveform_sig_rx =-1250;
32241: waveform_sig_rx =-1211;
32242: waveform_sig_rx =-930;
32243: waveform_sig_rx =-1197;
32244: waveform_sig_rx =-1219;
32245: waveform_sig_rx =-1070;
32246: waveform_sig_rx =-1035;
32247: waveform_sig_rx =-1307;
32248: waveform_sig_rx =-1075;
32249: waveform_sig_rx =-1044;
32250: waveform_sig_rx =-1246;
32251: waveform_sig_rx =-1190;
32252: waveform_sig_rx =-1006;
32253: waveform_sig_rx =-1132;
32254: waveform_sig_rx =-1315;
32255: waveform_sig_rx =-960;
32256: waveform_sig_rx =-1098;
32257: waveform_sig_rx =-1332;
32258: waveform_sig_rx =-1011;
32259: waveform_sig_rx =-1061;
32260: waveform_sig_rx =-1322;
32261: waveform_sig_rx =-1023;
32262: waveform_sig_rx =-1249;
32263: waveform_sig_rx =-1099;
32264: waveform_sig_rx =-1152;
32265: waveform_sig_rx =-1125;
32266: waveform_sig_rx =-1213;
32267: waveform_sig_rx =-1127;
32268: waveform_sig_rx =-1049;
32269: waveform_sig_rx =-1344;
32270: waveform_sig_rx =-1050;
32271: waveform_sig_rx =-1109;
32272: waveform_sig_rx =-1305;
32273: waveform_sig_rx =-1095;
32274: waveform_sig_rx =-1014;
32275: waveform_sig_rx =-1392;
32276: waveform_sig_rx =-1106;
32277: waveform_sig_rx =-997;
32278: waveform_sig_rx =-1404;
32279: waveform_sig_rx =-1098;
32280: waveform_sig_rx =-1026;
32281: waveform_sig_rx =-1287;
32282: waveform_sig_rx =-1215;
32283: waveform_sig_rx =-988;
32284: waveform_sig_rx =-1225;
32285: waveform_sig_rx =-1238;
32286: waveform_sig_rx =-1094;
32287: waveform_sig_rx =-1052;
32288: waveform_sig_rx =-1301;
32289: waveform_sig_rx =-1081;
32290: waveform_sig_rx =-1045;
32291: waveform_sig_rx =-1253;
32292: waveform_sig_rx =-1213;
32293: waveform_sig_rx =-974;
32294: waveform_sig_rx =-1167;
32295: waveform_sig_rx =-1331;
32296: waveform_sig_rx =-939;
32297: waveform_sig_rx =-1167;
32298: waveform_sig_rx =-1304;
32299: waveform_sig_rx =-979;
32300: waveform_sig_rx =-1089;
32301: waveform_sig_rx =-1259;
32302: waveform_sig_rx =-1041;
32303: waveform_sig_rx =-1270;
32304: waveform_sig_rx =-1032;
32305: waveform_sig_rx =-1197;
32306: waveform_sig_rx =-1065;
32307: waveform_sig_rx =-1192;
32308: waveform_sig_rx =-1188;
32309: waveform_sig_rx =-980;
32310: waveform_sig_rx =-1350;
32311: waveform_sig_rx =-1030;
32312: waveform_sig_rx =-1015;
32313: waveform_sig_rx =-1366;
32314: waveform_sig_rx =-981;
32315: waveform_sig_rx =-993;
32316: waveform_sig_rx =-1391;
32317: waveform_sig_rx =-978;
32318: waveform_sig_rx =-1007;
32319: waveform_sig_rx =-1336;
32320: waveform_sig_rx =-1022;
32321: waveform_sig_rx =-1007;
32322: waveform_sig_rx =-1232;
32323: waveform_sig_rx =-1155;
32324: waveform_sig_rx =-947;
32325: waveform_sig_rx =-1186;
32326: waveform_sig_rx =-1148;
32327: waveform_sig_rx =-1053;
32328: waveform_sig_rx =-982;
32329: waveform_sig_rx =-1246;
32330: waveform_sig_rx =-1074;
32331: waveform_sig_rx =-946;
32332: waveform_sig_rx =-1243;
32333: waveform_sig_rx =-1147;
32334: waveform_sig_rx =-890;
32335: waveform_sig_rx =-1204;
32336: waveform_sig_rx =-1166;
32337: waveform_sig_rx =-904;
32338: waveform_sig_rx =-1127;
32339: waveform_sig_rx =-1171;
32340: waveform_sig_rx =-992;
32341: waveform_sig_rx =-991;
32342: waveform_sig_rx =-1192;
32343: waveform_sig_rx =-1000;
32344: waveform_sig_rx =-1125;
32345: waveform_sig_rx =-974;
32346: waveform_sig_rx =-1130;
32347: waveform_sig_rx =-968;
32348: waveform_sig_rx =-1143;
32349: waveform_sig_rx =-1054;
32350: waveform_sig_rx =-868;
32351: waveform_sig_rx =-1295;
32352: waveform_sig_rx =-891;
32353: waveform_sig_rx =-948;
32354: waveform_sig_rx =-1278;
32355: waveform_sig_rx =-810;
32356: waveform_sig_rx =-949;
32357: waveform_sig_rx =-1261;
32358: waveform_sig_rx =-818;
32359: waveform_sig_rx =-961;
32360: waveform_sig_rx =-1161;
32361: waveform_sig_rx =-908;
32362: waveform_sig_rx =-911;
32363: waveform_sig_rx =-1078;
32364: waveform_sig_rx =-1058;
32365: waveform_sig_rx =-817;
32366: waveform_sig_rx =-1027;
32367: waveform_sig_rx =-1035;
32368: waveform_sig_rx =-891;
32369: waveform_sig_rx =-846;
32370: waveform_sig_rx =-1163;
32371: waveform_sig_rx =-880;
32372: waveform_sig_rx =-818;
32373: waveform_sig_rx =-1143;
32374: waveform_sig_rx =-936;
32375: waveform_sig_rx =-792;
32376: waveform_sig_rx =-1073;
32377: waveform_sig_rx =-996;
32378: waveform_sig_rx =-809;
32379: waveform_sig_rx =-939;
32380: waveform_sig_rx =-1049;
32381: waveform_sig_rx =-854;
32382: waveform_sig_rx =-804;
32383: waveform_sig_rx =-1085;
32384: waveform_sig_rx =-819;
32385: waveform_sig_rx =-963;
32386: waveform_sig_rx =-866;
32387: waveform_sig_rx =-937;
32388: waveform_sig_rx =-792;
32389: waveform_sig_rx =-1024;
32390: waveform_sig_rx =-817;
32391: waveform_sig_rx =-745;
32392: waveform_sig_rx =-1129;
32393: waveform_sig_rx =-649;
32394: waveform_sig_rx =-854;
32395: waveform_sig_rx =-1071;
32396: waveform_sig_rx =-642;
32397: waveform_sig_rx =-822;
32398: waveform_sig_rx =-1059;
32399: waveform_sig_rx =-660;
32400: waveform_sig_rx =-796;
32401: waveform_sig_rx =-946;
32402: waveform_sig_rx =-742;
32403: waveform_sig_rx =-736;
32404: waveform_sig_rx =-900;
32405: waveform_sig_rx =-882;
32406: waveform_sig_rx =-599;
32407: waveform_sig_rx =-875;
32408: waveform_sig_rx =-896;
32409: waveform_sig_rx =-673;
32410: waveform_sig_rx =-695;
32411: waveform_sig_rx =-962;
32412: waveform_sig_rx =-629;
32413: waveform_sig_rx =-687;
32414: waveform_sig_rx =-899;
32415: waveform_sig_rx =-712;
32416: waveform_sig_rx =-624;
32417: waveform_sig_rx =-803;
32418: waveform_sig_rx =-812;
32419: waveform_sig_rx =-598;
32420: waveform_sig_rx =-695;
32421: waveform_sig_rx =-877;
32422: waveform_sig_rx =-581;
32423: waveform_sig_rx =-592;
32424: waveform_sig_rx =-889;
32425: waveform_sig_rx =-521;
32426: waveform_sig_rx =-788;
32427: waveform_sig_rx =-616;
32428: waveform_sig_rx =-696;
32429: waveform_sig_rx =-609;
32430: waveform_sig_rx =-792;
32431: waveform_sig_rx =-560;
32432: waveform_sig_rx =-583;
32433: waveform_sig_rx =-848;
32434: waveform_sig_rx =-446;
32435: waveform_sig_rx =-653;
32436: waveform_sig_rx =-793;
32437: waveform_sig_rx =-430;
32438: waveform_sig_rx =-612;
32439: waveform_sig_rx =-783;
32440: waveform_sig_rx =-443;
32441: waveform_sig_rx =-554;
32442: waveform_sig_rx =-734;
32443: waveform_sig_rx =-536;
32444: waveform_sig_rx =-465;
32445: waveform_sig_rx =-688;
32446: waveform_sig_rx =-633;
32447: waveform_sig_rx =-338;
32448: waveform_sig_rx =-674;
32449: waveform_sig_rx =-615;
32450: waveform_sig_rx =-404;
32451: waveform_sig_rx =-491;
32452: waveform_sig_rx =-663;
32453: waveform_sig_rx =-393;
32454: waveform_sig_rx =-445;
32455: waveform_sig_rx =-594;
32456: waveform_sig_rx =-498;
32457: waveform_sig_rx =-343;
32458: waveform_sig_rx =-530;
32459: waveform_sig_rx =-598;
32460: waveform_sig_rx =-270;
32461: waveform_sig_rx =-483;
32462: waveform_sig_rx =-631;
32463: waveform_sig_rx =-260;
32464: waveform_sig_rx =-431;
32465: waveform_sig_rx =-589;
32466: waveform_sig_rx =-272;
32467: waveform_sig_rx =-569;
32468: waveform_sig_rx =-299;
32469: waveform_sig_rx =-479;
32470: waveform_sig_rx =-342;
32471: waveform_sig_rx =-502;
32472: waveform_sig_rx =-334;
32473: waveform_sig_rx =-323;
32474: waveform_sig_rx =-585;
32475: waveform_sig_rx =-180;
32476: waveform_sig_rx =-383;
32477: waveform_sig_rx =-515;
32478: waveform_sig_rx =-176;
32479: waveform_sig_rx =-333;
32480: waveform_sig_rx =-511;
32481: waveform_sig_rx =-200;
32482: waveform_sig_rx =-255;
32483: waveform_sig_rx =-470;
32484: waveform_sig_rx =-244;
32485: waveform_sig_rx =-155;
32486: waveform_sig_rx =-486;
32487: waveform_sig_rx =-303;
32488: waveform_sig_rx =-89;
32489: waveform_sig_rx =-432;
32490: waveform_sig_rx =-260;
32491: waveform_sig_rx =-200;
32492: waveform_sig_rx =-207;
32493: waveform_sig_rx =-363;
32494: waveform_sig_rx =-174;
32495: waveform_sig_rx =-116;
32496: waveform_sig_rx =-381;
32497: waveform_sig_rx =-212;
32498: waveform_sig_rx =-21;
32499: waveform_sig_rx =-326;
32500: waveform_sig_rx =-258;
32501: waveform_sig_rx =-10;
32502: waveform_sig_rx =-254;
32503: waveform_sig_rx =-304;
32504: waveform_sig_rx =10;
32505: waveform_sig_rx =-155;
32506: waveform_sig_rx =-273;
32507: waveform_sig_rx =-7;
32508: waveform_sig_rx =-276;
32509: waveform_sig_rx =5;
32510: waveform_sig_rx =-196;
32511: waveform_sig_rx =-32;
32512: waveform_sig_rx =-212;
32513: waveform_sig_rx =-30;
32514: waveform_sig_rx =-29;
32515: waveform_sig_rx =-276;
32516: waveform_sig_rx =77;
32517: waveform_sig_rx =-55;
32518: waveform_sig_rx =-251;
32519: waveform_sig_rx =128;
32520: waveform_sig_rx =-25;
32521: waveform_sig_rx =-281;
32522: waveform_sig_rx =175;
32523: waveform_sig_rx =-16;
32524: waveform_sig_rx =-205;
32525: waveform_sig_rx =118;
32526: waveform_sig_rx =65;
32527: waveform_sig_rx =-185;
32528: waveform_sig_rx =24;
32529: waveform_sig_rx =131;
32530: waveform_sig_rx =-80;
32531: waveform_sig_rx =1;
32532: waveform_sig_rx =110;
32533: waveform_sig_rx =117;
32534: waveform_sig_rx =-125;
32535: waveform_sig_rx =160;
32536: waveform_sig_rx =172;
32537: waveform_sig_rx =-108;
32538: waveform_sig_rx =109;
32539: waveform_sig_rx =262;
32540: waveform_sig_rx =-56;
32541: waveform_sig_rx =48;
32542: waveform_sig_rx =289;
32543: waveform_sig_rx =19;
32544: waveform_sig_rx =12;
32545: waveform_sig_rx =275;
32546: waveform_sig_rx =132;
32547: waveform_sig_rx =59;
32548: waveform_sig_rx =239;
32549: waveform_sig_rx =49;
32550: waveform_sig_rx =301;
32551: waveform_sig_rx =40;
32552: waveform_sig_rx =304;
32553: waveform_sig_rx =52;
32554: waveform_sig_rx =250;
32555: waveform_sig_rx =295;
32556: waveform_sig_rx =-29;
32557: waveform_sig_rx =425;
32558: waveform_sig_rx =233;
32559: waveform_sig_rx =5;
32560: waveform_sig_rx =521;
32561: waveform_sig_rx =212;
32562: waveform_sig_rx =43;
32563: waveform_sig_rx =489;
32564: waveform_sig_rx =229;
32565: waveform_sig_rx =134;
32566: waveform_sig_rx =414;
32567: waveform_sig_rx =357;
32568: waveform_sig_rx =143;
32569: waveform_sig_rx =334;
32570: waveform_sig_rx =443;
32571: waveform_sig_rx =225;
32572: waveform_sig_rx =264;
32573: waveform_sig_rx =406;
32574: waveform_sig_rx =382;
32575: waveform_sig_rx =149;
32576: waveform_sig_rx =479;
32577: waveform_sig_rx =433;
32578: waveform_sig_rx =164;
32579: waveform_sig_rx =441;
32580: waveform_sig_rx =518;
32581: waveform_sig_rx =223;
32582: waveform_sig_rx =395;
32583: waveform_sig_rx =538;
32584: waveform_sig_rx =307;
32585: waveform_sig_rx =326;
32586: waveform_sig_rx =524;
32587: waveform_sig_rx =467;
32588: waveform_sig_rx =323;
32589: waveform_sig_rx =509;
32590: waveform_sig_rx =403;
32591: waveform_sig_rx =499;
32592: waveform_sig_rx =379;
32593: waveform_sig_rx =587;
32594: waveform_sig_rx =268;
32595: waveform_sig_rx =621;
32596: waveform_sig_rx =497;
32597: waveform_sig_rx =283;
32598: waveform_sig_rx =749;
32599: waveform_sig_rx =414;
32600: waveform_sig_rx =352;
32601: waveform_sig_rx =749;
32602: waveform_sig_rx =462;
32603: waveform_sig_rx =339;
32604: waveform_sig_rx =762;
32605: waveform_sig_rx =495;
32606: waveform_sig_rx =397;
32607: waveform_sig_rx =688;
32608: waveform_sig_rx =589;
32609: waveform_sig_rx =437;
32610: waveform_sig_rx =569;
32611: waveform_sig_rx =683;
32612: waveform_sig_rx =530;
32613: waveform_sig_rx =462;
32614: waveform_sig_rx =747;
32615: waveform_sig_rx =614;
32616: waveform_sig_rx =363;
32617: waveform_sig_rx =831;
32618: waveform_sig_rx =600;
32619: waveform_sig_rx =483;
32620: waveform_sig_rx =725;
32621: waveform_sig_rx =726;
32622: waveform_sig_rx =568;
32623: waveform_sig_rx =594;
32624: waveform_sig_rx =816;
32625: waveform_sig_rx =603;
32626: waveform_sig_rx =546;
32627: waveform_sig_rx =843;
32628: waveform_sig_rx =683;
32629: waveform_sig_rx =571;
32630: waveform_sig_rx =774;
32631: waveform_sig_rx =620;
32632: waveform_sig_rx =757;
32633: waveform_sig_rx =648;
32634: waveform_sig_rx =822;
32635: waveform_sig_rx =519;
32636: waveform_sig_rx =912;
32637: waveform_sig_rx =702;
32638: waveform_sig_rx =551;
32639: waveform_sig_rx =979;
32640: waveform_sig_rx =609;
32641: waveform_sig_rx =636;
32642: waveform_sig_rx =975;
32643: waveform_sig_rx =651;
32644: waveform_sig_rx =635;
32645: waveform_sig_rx =956;
32646: waveform_sig_rx =733;
32647: waveform_sig_rx =680;
32648: waveform_sig_rx =864;
32649: waveform_sig_rx =852;
32650: waveform_sig_rx =661;
32651: waveform_sig_rx =795;
32652: waveform_sig_rx =976;
32653: waveform_sig_rx =701;
32654: waveform_sig_rx =734;
32655: waveform_sig_rx =1017;
32656: waveform_sig_rx =757;
32657: waveform_sig_rx =715;
32658: waveform_sig_rx =1025;
32659: waveform_sig_rx =795;
32660: waveform_sig_rx =773;
32661: waveform_sig_rx =884;
32662: waveform_sig_rx =989;
32663: waveform_sig_rx =748;
32664: waveform_sig_rx =800;
32665: waveform_sig_rx =1082;
32666: waveform_sig_rx =767;
32667: waveform_sig_rx =782;
32668: waveform_sig_rx =1076;
32669: waveform_sig_rx =858;
32670: waveform_sig_rx =803;
32671: waveform_sig_rx =981;
32672: waveform_sig_rx =819;
32673: waveform_sig_rx =970;
32674: waveform_sig_rx =884;
32675: waveform_sig_rx =994;
32676: waveform_sig_rx =737;
32677: waveform_sig_rx =1121;
32678: waveform_sig_rx =838;
32679: waveform_sig_rx =819;
32680: waveform_sig_rx =1143;
32681: waveform_sig_rx =776;
32682: waveform_sig_rx =903;
32683: waveform_sig_rx =1084;
32684: waveform_sig_rx =899;
32685: waveform_sig_rx =816;
32686: waveform_sig_rx =1113;
32687: waveform_sig_rx =969;
32688: waveform_sig_rx =799;
32689: waveform_sig_rx =1105;
32690: waveform_sig_rx =1061;
32691: waveform_sig_rx =750;
32692: waveform_sig_rx =1060;
32693: waveform_sig_rx =1114;
32694: waveform_sig_rx =861;
32695: waveform_sig_rx =982;
32696: waveform_sig_rx =1134;
32697: waveform_sig_rx =973;
32698: waveform_sig_rx =871;
32699: waveform_sig_rx =1163;
32700: waveform_sig_rx =993;
32701: waveform_sig_rx =892;
32702: waveform_sig_rx =1052;
32703: waveform_sig_rx =1146;
32704: waveform_sig_rx =874;
32705: waveform_sig_rx =954;
32706: waveform_sig_rx =1235;
32707: waveform_sig_rx =886;
32708: waveform_sig_rx =931;
32709: waveform_sig_rx =1257;
32710: waveform_sig_rx =942;
32711: waveform_sig_rx =986;
32712: waveform_sig_rx =1147;
32713: waveform_sig_rx =921;
32714: waveform_sig_rx =1169;
32715: waveform_sig_rx =975;
32716: waveform_sig_rx =1119;
32717: waveform_sig_rx =928;
32718: waveform_sig_rx =1232;
32719: waveform_sig_rx =1007;
32720: waveform_sig_rx =985;
32721: waveform_sig_rx =1227;
32722: waveform_sig_rx =1008;
32723: waveform_sig_rx =986;
32724: waveform_sig_rx =1259;
32725: waveform_sig_rx =1043;
32726: waveform_sig_rx =880;
32727: waveform_sig_rx =1341;
32728: waveform_sig_rx =1051;
32729: waveform_sig_rx =927;
32730: waveform_sig_rx =1285;
32731: waveform_sig_rx =1108;
32732: waveform_sig_rx =915;
32733: waveform_sig_rx =1204;
32734: waveform_sig_rx =1180;
32735: waveform_sig_rx =1007;
32736: waveform_sig_rx =1092;
32737: waveform_sig_rx =1237;
32738: waveform_sig_rx =1089;
32739: waveform_sig_rx =1012;
32740: waveform_sig_rx =1268;
32741: waveform_sig_rx =1154;
32742: waveform_sig_rx =1001;
32743: waveform_sig_rx =1175;
32744: waveform_sig_rx =1289;
32745: waveform_sig_rx =912;
32746: waveform_sig_rx =1141;
32747: waveform_sig_rx =1346;
32748: waveform_sig_rx =934;
32749: waveform_sig_rx =1121;
32750: waveform_sig_rx =1297;
32751: waveform_sig_rx =1018;
32752: waveform_sig_rx =1141;
32753: waveform_sig_rx =1137;
32754: waveform_sig_rx =1060;
32755: waveform_sig_rx =1252;
32756: waveform_sig_rx =996;
32757: waveform_sig_rx =1261;
32758: waveform_sig_rx =960;
32759: waveform_sig_rx =1288;
32760: waveform_sig_rx =1117;
32761: waveform_sig_rx =993;
32762: waveform_sig_rx =1345;
32763: waveform_sig_rx =1058;
32764: waveform_sig_rx =1006;
32765: waveform_sig_rx =1391;
32766: waveform_sig_rx =1037;
32767: waveform_sig_rx =995;


///////////////////////////////////////////////////

default: waveform_sig_rx= 0;
endcase

m_axis_src_data_tdata[15:0] = waveform_sig_rx;
m_axis_src_data_tdata[31:16] = waveform_sig_loopback; 



msg_count_tx_idx = msg_count_tx_idx + 1;
end else begin
m_axis_src_data_tvalid = 0;
end
end
endmodule
